magic
tech sky130A
magscale 1 2
timestamp 1762543975
<< viali >>
rect 17417 18785 17451 18819
rect 17509 18785 17543 18819
rect 16589 18717 16623 18751
rect 17785 18717 17819 18751
rect 18337 18717 18371 18751
rect 17325 18581 17359 18615
rect 17693 18581 17727 18615
rect 18061 18377 18095 18411
rect 16589 18241 16623 18275
rect 16313 18173 16347 18207
rect 18153 18173 18187 18207
rect 18245 18105 18279 18139
rect 19073 17765 19107 17799
rect 17601 17493 17635 17527
rect 16589 17153 16623 17187
rect 17969 17153 18003 17187
rect 18245 17085 18279 17119
rect 14105 16745 14139 16779
rect 18613 16745 18647 16779
rect 15393 16677 15427 16711
rect 17325 16677 17359 16711
rect 19073 9877 19107 9911
rect 3801 765 3835 799
rect 6285 765 6319 799
rect 8769 765 8803 799
rect 11253 765 11287 799
rect 13737 765 13771 799
rect 16221 765 16255 799
rect 18705 765 18739 799
<< metal1 >>
rect 552 19066 19571 19088
rect 552 19014 5112 19066
rect 5164 19014 5176 19066
rect 5228 19014 5240 19066
rect 5292 19014 5304 19066
rect 5356 19014 5368 19066
rect 5420 19014 9827 19066
rect 9879 19014 9891 19066
rect 9943 19014 9955 19066
rect 10007 19014 10019 19066
rect 10071 19014 10083 19066
rect 10135 19014 14542 19066
rect 14594 19014 14606 19066
rect 14658 19014 14670 19066
rect 14722 19014 14734 19066
rect 14786 19014 14798 19066
rect 14850 19014 19257 19066
rect 19309 19014 19321 19066
rect 19373 19014 19385 19066
rect 19437 19014 19449 19066
rect 19501 19014 19513 19066
rect 19565 19014 19571 19066
rect 552 18992 19571 19014
rect 17402 18912 17408 18964
rect 17460 18912 17466 18964
rect 17420 18884 17448 18912
rect 17420 18856 17540 18884
rect 17512 18825 17540 18856
rect 17405 18819 17463 18825
rect 17405 18785 17417 18819
rect 17451 18785 17463 18819
rect 17405 18779 17463 18785
rect 17497 18819 17555 18825
rect 17497 18785 17509 18819
rect 17543 18785 17555 18819
rect 17497 18779 17555 18785
rect 16574 18708 16580 18760
rect 16632 18708 16638 18760
rect 17420 18748 17448 18779
rect 17773 18751 17831 18757
rect 17773 18748 17785 18751
rect 17420 18720 17785 18748
rect 17773 18717 17785 18720
rect 17819 18717 17831 18751
rect 17773 18711 17831 18717
rect 18322 18708 18328 18760
rect 18380 18708 18386 18760
rect 17310 18572 17316 18624
rect 17368 18572 17374 18624
rect 17678 18572 17684 18624
rect 17736 18572 17742 18624
rect 552 18522 19412 18544
rect 552 18470 2755 18522
rect 2807 18470 2819 18522
rect 2871 18470 2883 18522
rect 2935 18470 2947 18522
rect 2999 18470 3011 18522
rect 3063 18470 7470 18522
rect 7522 18470 7534 18522
rect 7586 18470 7598 18522
rect 7650 18470 7662 18522
rect 7714 18470 7726 18522
rect 7778 18470 12185 18522
rect 12237 18470 12249 18522
rect 12301 18470 12313 18522
rect 12365 18470 12377 18522
rect 12429 18470 12441 18522
rect 12493 18470 16900 18522
rect 16952 18470 16964 18522
rect 17016 18470 17028 18522
rect 17080 18470 17092 18522
rect 17144 18470 17156 18522
rect 17208 18470 19412 18522
rect 552 18448 19412 18470
rect 17678 18368 17684 18420
rect 17736 18368 17742 18420
rect 18049 18411 18107 18417
rect 18049 18377 18061 18411
rect 18095 18408 18107 18411
rect 18322 18408 18328 18420
rect 18095 18380 18328 18408
rect 18095 18377 18107 18380
rect 18049 18371 18107 18377
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 16574 18232 16580 18284
rect 16632 18232 16638 18284
rect 17696 18272 17724 18368
rect 17696 18244 18184 18272
rect 14090 18164 14096 18216
rect 14148 18204 14154 18216
rect 18156 18213 18184 18244
rect 16301 18207 16359 18213
rect 16301 18204 16313 18207
rect 14148 18176 16313 18204
rect 14148 18164 14154 18176
rect 16301 18173 16313 18176
rect 16347 18173 16359 18207
rect 16301 18167 16359 18173
rect 18141 18207 18199 18213
rect 18141 18173 18153 18207
rect 18187 18173 18199 18207
rect 18141 18167 18199 18173
rect 18233 18139 18291 18145
rect 18233 18136 18245 18139
rect 17802 18108 18245 18136
rect 18233 18105 18245 18108
rect 18279 18105 18291 18139
rect 18233 18099 18291 18105
rect 552 17978 19571 18000
rect 552 17926 5112 17978
rect 5164 17926 5176 17978
rect 5228 17926 5240 17978
rect 5292 17926 5304 17978
rect 5356 17926 5368 17978
rect 5420 17926 9827 17978
rect 9879 17926 9891 17978
rect 9943 17926 9955 17978
rect 10007 17926 10019 17978
rect 10071 17926 10083 17978
rect 10135 17926 14542 17978
rect 14594 17926 14606 17978
rect 14658 17926 14670 17978
rect 14722 17926 14734 17978
rect 14786 17926 14798 17978
rect 14850 17926 19257 17978
rect 19309 17926 19321 17978
rect 19373 17926 19385 17978
rect 19437 17926 19449 17978
rect 19501 17926 19513 17978
rect 19565 17926 19571 17978
rect 552 17904 19571 17926
rect 19058 17756 19064 17808
rect 19116 17756 19122 17808
rect 17586 17484 17592 17536
rect 17644 17484 17650 17536
rect 552 17434 19412 17456
rect 552 17382 2755 17434
rect 2807 17382 2819 17434
rect 2871 17382 2883 17434
rect 2935 17382 2947 17434
rect 2999 17382 3011 17434
rect 3063 17382 7470 17434
rect 7522 17382 7534 17434
rect 7586 17382 7598 17434
rect 7650 17382 7662 17434
rect 7714 17382 7726 17434
rect 7778 17382 12185 17434
rect 12237 17382 12249 17434
rect 12301 17382 12313 17434
rect 12365 17382 12377 17434
rect 12429 17382 12441 17434
rect 12493 17382 16900 17434
rect 16952 17382 16964 17434
rect 17016 17382 17028 17434
rect 17080 17382 17092 17434
rect 17144 17382 17156 17434
rect 17208 17382 19412 17434
rect 552 17360 19412 17382
rect 1210 17212 1216 17264
rect 1268 17252 1274 17264
rect 1268 17224 9674 17252
rect 1268 17212 1274 17224
rect 9646 17184 9674 17224
rect 16577 17187 16635 17193
rect 16577 17184 16589 17187
rect 9646 17156 16589 17184
rect 16577 17153 16589 17156
rect 16623 17153 16635 17187
rect 16577 17147 16635 17153
rect 17310 17144 17316 17196
rect 17368 17184 17374 17196
rect 17957 17187 18015 17193
rect 17957 17184 17969 17187
rect 17368 17156 17969 17184
rect 17368 17144 17374 17156
rect 17957 17153 17969 17156
rect 18003 17153 18015 17187
rect 17957 17147 18015 17153
rect 18233 17119 18291 17125
rect 18233 17085 18245 17119
rect 18279 17116 18291 17119
rect 18598 17116 18604 17128
rect 18279 17088 18604 17116
rect 18279 17085 18291 17088
rect 18233 17079 18291 17085
rect 18598 17076 18604 17088
rect 18656 17076 18662 17128
rect 552 16890 19571 16912
rect 552 16838 5112 16890
rect 5164 16838 5176 16890
rect 5228 16838 5240 16890
rect 5292 16838 5304 16890
rect 5356 16838 5368 16890
rect 5420 16838 9827 16890
rect 9879 16838 9891 16890
rect 9943 16838 9955 16890
rect 10007 16838 10019 16890
rect 10071 16838 10083 16890
rect 10135 16838 14542 16890
rect 14594 16838 14606 16890
rect 14658 16838 14670 16890
rect 14722 16838 14734 16890
rect 14786 16838 14798 16890
rect 14850 16838 19257 16890
rect 19309 16838 19321 16890
rect 19373 16838 19385 16890
rect 19437 16838 19449 16890
rect 19501 16838 19513 16890
rect 19565 16838 19571 16890
rect 552 16816 19571 16838
rect 14090 16736 14096 16788
rect 14148 16736 14154 16788
rect 17586 16736 17592 16788
rect 17644 16736 17650 16788
rect 18598 16736 18604 16788
rect 18656 16736 18662 16788
rect 15381 16711 15439 16717
rect 15381 16677 15393 16711
rect 15427 16708 15439 16711
rect 17313 16711 17371 16717
rect 17313 16708 17325 16711
rect 15427 16680 17325 16708
rect 15427 16677 15439 16680
rect 15381 16671 15439 16677
rect 17313 16677 17325 16680
rect 17359 16708 17371 16711
rect 17604 16708 17632 16736
rect 17359 16680 17632 16708
rect 17359 16677 17371 16680
rect 17313 16671 17371 16677
rect 552 16346 19412 16368
rect 552 16294 2755 16346
rect 2807 16294 2819 16346
rect 2871 16294 2883 16346
rect 2935 16294 2947 16346
rect 2999 16294 3011 16346
rect 3063 16294 7470 16346
rect 7522 16294 7534 16346
rect 7586 16294 7598 16346
rect 7650 16294 7662 16346
rect 7714 16294 7726 16346
rect 7778 16294 12185 16346
rect 12237 16294 12249 16346
rect 12301 16294 12313 16346
rect 12365 16294 12377 16346
rect 12429 16294 12441 16346
rect 12493 16294 16900 16346
rect 16952 16294 16964 16346
rect 17016 16294 17028 16346
rect 17080 16294 17092 16346
rect 17144 16294 17156 16346
rect 17208 16294 19412 16346
rect 552 16272 19412 16294
rect 552 15802 19571 15824
rect 552 15750 5112 15802
rect 5164 15750 5176 15802
rect 5228 15750 5240 15802
rect 5292 15750 5304 15802
rect 5356 15750 5368 15802
rect 5420 15750 9827 15802
rect 9879 15750 9891 15802
rect 9943 15750 9955 15802
rect 10007 15750 10019 15802
rect 10071 15750 10083 15802
rect 10135 15750 14542 15802
rect 14594 15750 14606 15802
rect 14658 15750 14670 15802
rect 14722 15750 14734 15802
rect 14786 15750 14798 15802
rect 14850 15750 19257 15802
rect 19309 15750 19321 15802
rect 19373 15750 19385 15802
rect 19437 15750 19449 15802
rect 19501 15750 19513 15802
rect 19565 15750 19571 15802
rect 552 15728 19571 15750
rect 552 15258 19412 15280
rect 552 15206 2755 15258
rect 2807 15206 2819 15258
rect 2871 15206 2883 15258
rect 2935 15206 2947 15258
rect 2999 15206 3011 15258
rect 3063 15206 7470 15258
rect 7522 15206 7534 15258
rect 7586 15206 7598 15258
rect 7650 15206 7662 15258
rect 7714 15206 7726 15258
rect 7778 15206 12185 15258
rect 12237 15206 12249 15258
rect 12301 15206 12313 15258
rect 12365 15206 12377 15258
rect 12429 15206 12441 15258
rect 12493 15206 16900 15258
rect 16952 15206 16964 15258
rect 17016 15206 17028 15258
rect 17080 15206 17092 15258
rect 17144 15206 17156 15258
rect 17208 15206 19412 15258
rect 552 15184 19412 15206
rect 552 14714 19571 14736
rect 552 14662 5112 14714
rect 5164 14662 5176 14714
rect 5228 14662 5240 14714
rect 5292 14662 5304 14714
rect 5356 14662 5368 14714
rect 5420 14662 9827 14714
rect 9879 14662 9891 14714
rect 9943 14662 9955 14714
rect 10007 14662 10019 14714
rect 10071 14662 10083 14714
rect 10135 14662 14542 14714
rect 14594 14662 14606 14714
rect 14658 14662 14670 14714
rect 14722 14662 14734 14714
rect 14786 14662 14798 14714
rect 14850 14662 19257 14714
rect 19309 14662 19321 14714
rect 19373 14662 19385 14714
rect 19437 14662 19449 14714
rect 19501 14662 19513 14714
rect 19565 14662 19571 14714
rect 552 14640 19571 14662
rect 552 14170 19412 14192
rect 552 14118 2755 14170
rect 2807 14118 2819 14170
rect 2871 14118 2883 14170
rect 2935 14118 2947 14170
rect 2999 14118 3011 14170
rect 3063 14118 7470 14170
rect 7522 14118 7534 14170
rect 7586 14118 7598 14170
rect 7650 14118 7662 14170
rect 7714 14118 7726 14170
rect 7778 14118 12185 14170
rect 12237 14118 12249 14170
rect 12301 14118 12313 14170
rect 12365 14118 12377 14170
rect 12429 14118 12441 14170
rect 12493 14118 16900 14170
rect 16952 14118 16964 14170
rect 17016 14118 17028 14170
rect 17080 14118 17092 14170
rect 17144 14118 17156 14170
rect 17208 14118 19412 14170
rect 552 14096 19412 14118
rect 552 13626 19571 13648
rect 552 13574 5112 13626
rect 5164 13574 5176 13626
rect 5228 13574 5240 13626
rect 5292 13574 5304 13626
rect 5356 13574 5368 13626
rect 5420 13574 9827 13626
rect 9879 13574 9891 13626
rect 9943 13574 9955 13626
rect 10007 13574 10019 13626
rect 10071 13574 10083 13626
rect 10135 13574 14542 13626
rect 14594 13574 14606 13626
rect 14658 13574 14670 13626
rect 14722 13574 14734 13626
rect 14786 13574 14798 13626
rect 14850 13574 19257 13626
rect 19309 13574 19321 13626
rect 19373 13574 19385 13626
rect 19437 13574 19449 13626
rect 19501 13574 19513 13626
rect 19565 13574 19571 13626
rect 552 13552 19571 13574
rect 552 13082 19412 13104
rect 552 13030 2755 13082
rect 2807 13030 2819 13082
rect 2871 13030 2883 13082
rect 2935 13030 2947 13082
rect 2999 13030 3011 13082
rect 3063 13030 7470 13082
rect 7522 13030 7534 13082
rect 7586 13030 7598 13082
rect 7650 13030 7662 13082
rect 7714 13030 7726 13082
rect 7778 13030 12185 13082
rect 12237 13030 12249 13082
rect 12301 13030 12313 13082
rect 12365 13030 12377 13082
rect 12429 13030 12441 13082
rect 12493 13030 16900 13082
rect 16952 13030 16964 13082
rect 17016 13030 17028 13082
rect 17080 13030 17092 13082
rect 17144 13030 17156 13082
rect 17208 13030 19412 13082
rect 552 13008 19412 13030
rect 552 12538 19571 12560
rect 552 12486 5112 12538
rect 5164 12486 5176 12538
rect 5228 12486 5240 12538
rect 5292 12486 5304 12538
rect 5356 12486 5368 12538
rect 5420 12486 9827 12538
rect 9879 12486 9891 12538
rect 9943 12486 9955 12538
rect 10007 12486 10019 12538
rect 10071 12486 10083 12538
rect 10135 12486 14542 12538
rect 14594 12486 14606 12538
rect 14658 12486 14670 12538
rect 14722 12486 14734 12538
rect 14786 12486 14798 12538
rect 14850 12486 19257 12538
rect 19309 12486 19321 12538
rect 19373 12486 19385 12538
rect 19437 12486 19449 12538
rect 19501 12486 19513 12538
rect 19565 12486 19571 12538
rect 552 12464 19571 12486
rect 552 11994 19412 12016
rect 552 11942 2755 11994
rect 2807 11942 2819 11994
rect 2871 11942 2883 11994
rect 2935 11942 2947 11994
rect 2999 11942 3011 11994
rect 3063 11942 7470 11994
rect 7522 11942 7534 11994
rect 7586 11942 7598 11994
rect 7650 11942 7662 11994
rect 7714 11942 7726 11994
rect 7778 11942 12185 11994
rect 12237 11942 12249 11994
rect 12301 11942 12313 11994
rect 12365 11942 12377 11994
rect 12429 11942 12441 11994
rect 12493 11942 16900 11994
rect 16952 11942 16964 11994
rect 17016 11942 17028 11994
rect 17080 11942 17092 11994
rect 17144 11942 17156 11994
rect 17208 11942 19412 11994
rect 552 11920 19412 11942
rect 552 11450 19571 11472
rect 552 11398 5112 11450
rect 5164 11398 5176 11450
rect 5228 11398 5240 11450
rect 5292 11398 5304 11450
rect 5356 11398 5368 11450
rect 5420 11398 9827 11450
rect 9879 11398 9891 11450
rect 9943 11398 9955 11450
rect 10007 11398 10019 11450
rect 10071 11398 10083 11450
rect 10135 11398 14542 11450
rect 14594 11398 14606 11450
rect 14658 11398 14670 11450
rect 14722 11398 14734 11450
rect 14786 11398 14798 11450
rect 14850 11398 19257 11450
rect 19309 11398 19321 11450
rect 19373 11398 19385 11450
rect 19437 11398 19449 11450
rect 19501 11398 19513 11450
rect 19565 11398 19571 11450
rect 552 11376 19571 11398
rect 552 10906 19412 10928
rect 552 10854 2755 10906
rect 2807 10854 2819 10906
rect 2871 10854 2883 10906
rect 2935 10854 2947 10906
rect 2999 10854 3011 10906
rect 3063 10854 7470 10906
rect 7522 10854 7534 10906
rect 7586 10854 7598 10906
rect 7650 10854 7662 10906
rect 7714 10854 7726 10906
rect 7778 10854 12185 10906
rect 12237 10854 12249 10906
rect 12301 10854 12313 10906
rect 12365 10854 12377 10906
rect 12429 10854 12441 10906
rect 12493 10854 16900 10906
rect 16952 10854 16964 10906
rect 17016 10854 17028 10906
rect 17080 10854 17092 10906
rect 17144 10854 17156 10906
rect 17208 10854 19412 10906
rect 552 10832 19412 10854
rect 552 10362 19571 10384
rect 552 10310 5112 10362
rect 5164 10310 5176 10362
rect 5228 10310 5240 10362
rect 5292 10310 5304 10362
rect 5356 10310 5368 10362
rect 5420 10310 9827 10362
rect 9879 10310 9891 10362
rect 9943 10310 9955 10362
rect 10007 10310 10019 10362
rect 10071 10310 10083 10362
rect 10135 10310 14542 10362
rect 14594 10310 14606 10362
rect 14658 10310 14670 10362
rect 14722 10310 14734 10362
rect 14786 10310 14798 10362
rect 14850 10310 19257 10362
rect 19309 10310 19321 10362
rect 19373 10310 19385 10362
rect 19437 10310 19449 10362
rect 19501 10310 19513 10362
rect 19565 10310 19571 10362
rect 552 10288 19571 10310
rect 19058 9868 19064 9920
rect 19116 9868 19122 9920
rect 552 9818 19412 9840
rect 552 9766 2755 9818
rect 2807 9766 2819 9818
rect 2871 9766 2883 9818
rect 2935 9766 2947 9818
rect 2999 9766 3011 9818
rect 3063 9766 7470 9818
rect 7522 9766 7534 9818
rect 7586 9766 7598 9818
rect 7650 9766 7662 9818
rect 7714 9766 7726 9818
rect 7778 9766 12185 9818
rect 12237 9766 12249 9818
rect 12301 9766 12313 9818
rect 12365 9766 12377 9818
rect 12429 9766 12441 9818
rect 12493 9766 16900 9818
rect 16952 9766 16964 9818
rect 17016 9766 17028 9818
rect 17080 9766 17092 9818
rect 17144 9766 17156 9818
rect 17208 9766 19412 9818
rect 552 9744 19412 9766
rect 552 9274 19571 9296
rect 552 9222 5112 9274
rect 5164 9222 5176 9274
rect 5228 9222 5240 9274
rect 5292 9222 5304 9274
rect 5356 9222 5368 9274
rect 5420 9222 9827 9274
rect 9879 9222 9891 9274
rect 9943 9222 9955 9274
rect 10007 9222 10019 9274
rect 10071 9222 10083 9274
rect 10135 9222 14542 9274
rect 14594 9222 14606 9274
rect 14658 9222 14670 9274
rect 14722 9222 14734 9274
rect 14786 9222 14798 9274
rect 14850 9222 19257 9274
rect 19309 9222 19321 9274
rect 19373 9222 19385 9274
rect 19437 9222 19449 9274
rect 19501 9222 19513 9274
rect 19565 9222 19571 9274
rect 552 9200 19571 9222
rect 552 8730 19412 8752
rect 552 8678 2755 8730
rect 2807 8678 2819 8730
rect 2871 8678 2883 8730
rect 2935 8678 2947 8730
rect 2999 8678 3011 8730
rect 3063 8678 7470 8730
rect 7522 8678 7534 8730
rect 7586 8678 7598 8730
rect 7650 8678 7662 8730
rect 7714 8678 7726 8730
rect 7778 8678 12185 8730
rect 12237 8678 12249 8730
rect 12301 8678 12313 8730
rect 12365 8678 12377 8730
rect 12429 8678 12441 8730
rect 12493 8678 16900 8730
rect 16952 8678 16964 8730
rect 17016 8678 17028 8730
rect 17080 8678 17092 8730
rect 17144 8678 17156 8730
rect 17208 8678 19412 8730
rect 552 8656 19412 8678
rect 552 8186 19571 8208
rect 552 8134 5112 8186
rect 5164 8134 5176 8186
rect 5228 8134 5240 8186
rect 5292 8134 5304 8186
rect 5356 8134 5368 8186
rect 5420 8134 9827 8186
rect 9879 8134 9891 8186
rect 9943 8134 9955 8186
rect 10007 8134 10019 8186
rect 10071 8134 10083 8186
rect 10135 8134 14542 8186
rect 14594 8134 14606 8186
rect 14658 8134 14670 8186
rect 14722 8134 14734 8186
rect 14786 8134 14798 8186
rect 14850 8134 19257 8186
rect 19309 8134 19321 8186
rect 19373 8134 19385 8186
rect 19437 8134 19449 8186
rect 19501 8134 19513 8186
rect 19565 8134 19571 8186
rect 552 8112 19571 8134
rect 552 7642 19412 7664
rect 552 7590 2755 7642
rect 2807 7590 2819 7642
rect 2871 7590 2883 7642
rect 2935 7590 2947 7642
rect 2999 7590 3011 7642
rect 3063 7590 7470 7642
rect 7522 7590 7534 7642
rect 7586 7590 7598 7642
rect 7650 7590 7662 7642
rect 7714 7590 7726 7642
rect 7778 7590 12185 7642
rect 12237 7590 12249 7642
rect 12301 7590 12313 7642
rect 12365 7590 12377 7642
rect 12429 7590 12441 7642
rect 12493 7590 16900 7642
rect 16952 7590 16964 7642
rect 17016 7590 17028 7642
rect 17080 7590 17092 7642
rect 17144 7590 17156 7642
rect 17208 7590 19412 7642
rect 552 7568 19412 7590
rect 552 7098 19571 7120
rect 552 7046 5112 7098
rect 5164 7046 5176 7098
rect 5228 7046 5240 7098
rect 5292 7046 5304 7098
rect 5356 7046 5368 7098
rect 5420 7046 9827 7098
rect 9879 7046 9891 7098
rect 9943 7046 9955 7098
rect 10007 7046 10019 7098
rect 10071 7046 10083 7098
rect 10135 7046 14542 7098
rect 14594 7046 14606 7098
rect 14658 7046 14670 7098
rect 14722 7046 14734 7098
rect 14786 7046 14798 7098
rect 14850 7046 19257 7098
rect 19309 7046 19321 7098
rect 19373 7046 19385 7098
rect 19437 7046 19449 7098
rect 19501 7046 19513 7098
rect 19565 7046 19571 7098
rect 552 7024 19571 7046
rect 552 6554 19412 6576
rect 552 6502 2755 6554
rect 2807 6502 2819 6554
rect 2871 6502 2883 6554
rect 2935 6502 2947 6554
rect 2999 6502 3011 6554
rect 3063 6502 7470 6554
rect 7522 6502 7534 6554
rect 7586 6502 7598 6554
rect 7650 6502 7662 6554
rect 7714 6502 7726 6554
rect 7778 6502 12185 6554
rect 12237 6502 12249 6554
rect 12301 6502 12313 6554
rect 12365 6502 12377 6554
rect 12429 6502 12441 6554
rect 12493 6502 16900 6554
rect 16952 6502 16964 6554
rect 17016 6502 17028 6554
rect 17080 6502 17092 6554
rect 17144 6502 17156 6554
rect 17208 6502 19412 6554
rect 552 6480 19412 6502
rect 552 6010 19571 6032
rect 552 5958 5112 6010
rect 5164 5958 5176 6010
rect 5228 5958 5240 6010
rect 5292 5958 5304 6010
rect 5356 5958 5368 6010
rect 5420 5958 9827 6010
rect 9879 5958 9891 6010
rect 9943 5958 9955 6010
rect 10007 5958 10019 6010
rect 10071 5958 10083 6010
rect 10135 5958 14542 6010
rect 14594 5958 14606 6010
rect 14658 5958 14670 6010
rect 14722 5958 14734 6010
rect 14786 5958 14798 6010
rect 14850 5958 19257 6010
rect 19309 5958 19321 6010
rect 19373 5958 19385 6010
rect 19437 5958 19449 6010
rect 19501 5958 19513 6010
rect 19565 5958 19571 6010
rect 552 5936 19571 5958
rect 552 5466 19412 5488
rect 552 5414 2755 5466
rect 2807 5414 2819 5466
rect 2871 5414 2883 5466
rect 2935 5414 2947 5466
rect 2999 5414 3011 5466
rect 3063 5414 7470 5466
rect 7522 5414 7534 5466
rect 7586 5414 7598 5466
rect 7650 5414 7662 5466
rect 7714 5414 7726 5466
rect 7778 5414 12185 5466
rect 12237 5414 12249 5466
rect 12301 5414 12313 5466
rect 12365 5414 12377 5466
rect 12429 5414 12441 5466
rect 12493 5414 16900 5466
rect 16952 5414 16964 5466
rect 17016 5414 17028 5466
rect 17080 5414 17092 5466
rect 17144 5414 17156 5466
rect 17208 5414 19412 5466
rect 552 5392 19412 5414
rect 552 4922 19571 4944
rect 552 4870 5112 4922
rect 5164 4870 5176 4922
rect 5228 4870 5240 4922
rect 5292 4870 5304 4922
rect 5356 4870 5368 4922
rect 5420 4870 9827 4922
rect 9879 4870 9891 4922
rect 9943 4870 9955 4922
rect 10007 4870 10019 4922
rect 10071 4870 10083 4922
rect 10135 4870 14542 4922
rect 14594 4870 14606 4922
rect 14658 4870 14670 4922
rect 14722 4870 14734 4922
rect 14786 4870 14798 4922
rect 14850 4870 19257 4922
rect 19309 4870 19321 4922
rect 19373 4870 19385 4922
rect 19437 4870 19449 4922
rect 19501 4870 19513 4922
rect 19565 4870 19571 4922
rect 552 4848 19571 4870
rect 552 4378 19412 4400
rect 552 4326 2755 4378
rect 2807 4326 2819 4378
rect 2871 4326 2883 4378
rect 2935 4326 2947 4378
rect 2999 4326 3011 4378
rect 3063 4326 7470 4378
rect 7522 4326 7534 4378
rect 7586 4326 7598 4378
rect 7650 4326 7662 4378
rect 7714 4326 7726 4378
rect 7778 4326 12185 4378
rect 12237 4326 12249 4378
rect 12301 4326 12313 4378
rect 12365 4326 12377 4378
rect 12429 4326 12441 4378
rect 12493 4326 16900 4378
rect 16952 4326 16964 4378
rect 17016 4326 17028 4378
rect 17080 4326 17092 4378
rect 17144 4326 17156 4378
rect 17208 4326 19412 4378
rect 552 4304 19412 4326
rect 552 3834 19571 3856
rect 552 3782 5112 3834
rect 5164 3782 5176 3834
rect 5228 3782 5240 3834
rect 5292 3782 5304 3834
rect 5356 3782 5368 3834
rect 5420 3782 9827 3834
rect 9879 3782 9891 3834
rect 9943 3782 9955 3834
rect 10007 3782 10019 3834
rect 10071 3782 10083 3834
rect 10135 3782 14542 3834
rect 14594 3782 14606 3834
rect 14658 3782 14670 3834
rect 14722 3782 14734 3834
rect 14786 3782 14798 3834
rect 14850 3782 19257 3834
rect 19309 3782 19321 3834
rect 19373 3782 19385 3834
rect 19437 3782 19449 3834
rect 19501 3782 19513 3834
rect 19565 3782 19571 3834
rect 552 3760 19571 3782
rect 552 3290 19412 3312
rect 552 3238 2755 3290
rect 2807 3238 2819 3290
rect 2871 3238 2883 3290
rect 2935 3238 2947 3290
rect 2999 3238 3011 3290
rect 3063 3238 7470 3290
rect 7522 3238 7534 3290
rect 7586 3238 7598 3290
rect 7650 3238 7662 3290
rect 7714 3238 7726 3290
rect 7778 3238 12185 3290
rect 12237 3238 12249 3290
rect 12301 3238 12313 3290
rect 12365 3238 12377 3290
rect 12429 3238 12441 3290
rect 12493 3238 16900 3290
rect 16952 3238 16964 3290
rect 17016 3238 17028 3290
rect 17080 3238 17092 3290
rect 17144 3238 17156 3290
rect 17208 3238 19412 3290
rect 552 3216 19412 3238
rect 552 2746 19571 2768
rect 552 2694 5112 2746
rect 5164 2694 5176 2746
rect 5228 2694 5240 2746
rect 5292 2694 5304 2746
rect 5356 2694 5368 2746
rect 5420 2694 9827 2746
rect 9879 2694 9891 2746
rect 9943 2694 9955 2746
rect 10007 2694 10019 2746
rect 10071 2694 10083 2746
rect 10135 2694 14542 2746
rect 14594 2694 14606 2746
rect 14658 2694 14670 2746
rect 14722 2694 14734 2746
rect 14786 2694 14798 2746
rect 14850 2694 19257 2746
rect 19309 2694 19321 2746
rect 19373 2694 19385 2746
rect 19437 2694 19449 2746
rect 19501 2694 19513 2746
rect 19565 2694 19571 2746
rect 552 2672 19571 2694
rect 552 2202 19412 2224
rect 552 2150 2755 2202
rect 2807 2150 2819 2202
rect 2871 2150 2883 2202
rect 2935 2150 2947 2202
rect 2999 2150 3011 2202
rect 3063 2150 7470 2202
rect 7522 2150 7534 2202
rect 7586 2150 7598 2202
rect 7650 2150 7662 2202
rect 7714 2150 7726 2202
rect 7778 2150 12185 2202
rect 12237 2150 12249 2202
rect 12301 2150 12313 2202
rect 12365 2150 12377 2202
rect 12429 2150 12441 2202
rect 12493 2150 16900 2202
rect 16952 2150 16964 2202
rect 17016 2150 17028 2202
rect 17080 2150 17092 2202
rect 17144 2150 17156 2202
rect 17208 2150 19412 2202
rect 552 2128 19412 2150
rect 552 1658 19571 1680
rect 552 1606 5112 1658
rect 5164 1606 5176 1658
rect 5228 1606 5240 1658
rect 5292 1606 5304 1658
rect 5356 1606 5368 1658
rect 5420 1606 9827 1658
rect 9879 1606 9891 1658
rect 9943 1606 9955 1658
rect 10007 1606 10019 1658
rect 10071 1606 10083 1658
rect 10135 1606 14542 1658
rect 14594 1606 14606 1658
rect 14658 1606 14670 1658
rect 14722 1606 14734 1658
rect 14786 1606 14798 1658
rect 14850 1606 19257 1658
rect 19309 1606 19321 1658
rect 19373 1606 19385 1658
rect 19437 1606 19449 1658
rect 19501 1606 19513 1658
rect 19565 1606 19571 1658
rect 552 1584 19571 1606
rect 552 1114 19412 1136
rect 552 1062 2755 1114
rect 2807 1062 2819 1114
rect 2871 1062 2883 1114
rect 2935 1062 2947 1114
rect 2999 1062 3011 1114
rect 3063 1062 7470 1114
rect 7522 1062 7534 1114
rect 7586 1062 7598 1114
rect 7650 1062 7662 1114
rect 7714 1062 7726 1114
rect 7778 1062 12185 1114
rect 12237 1062 12249 1114
rect 12301 1062 12313 1114
rect 12365 1062 12377 1114
rect 12429 1062 12441 1114
rect 12493 1062 16900 1114
rect 16952 1062 16964 1114
rect 17016 1062 17028 1114
rect 17080 1062 17092 1114
rect 17144 1062 17156 1114
rect 17208 1062 19412 1114
rect 552 1040 19412 1062
rect 3786 756 3792 808
rect 3844 756 3850 808
rect 6270 756 6276 808
rect 6328 756 6334 808
rect 8754 756 8760 808
rect 8812 756 8818 808
rect 11238 756 11244 808
rect 11296 756 11302 808
rect 13722 756 13728 808
rect 13780 756 13786 808
rect 16206 756 16212 808
rect 16264 756 16270 808
rect 18690 756 18696 808
rect 18748 756 18754 808
rect 552 570 19571 592
rect 552 518 5112 570
rect 5164 518 5176 570
rect 5228 518 5240 570
rect 5292 518 5304 570
rect 5356 518 5368 570
rect 5420 518 9827 570
rect 9879 518 9891 570
rect 9943 518 9955 570
rect 10007 518 10019 570
rect 10071 518 10083 570
rect 10135 518 14542 570
rect 14594 518 14606 570
rect 14658 518 14670 570
rect 14722 518 14734 570
rect 14786 518 14798 570
rect 14850 518 19257 570
rect 19309 518 19321 570
rect 19373 518 19385 570
rect 19437 518 19449 570
rect 19501 518 19513 570
rect 19565 518 19571 570
rect 552 496 19571 518
<< via1 >>
rect 5112 19014 5164 19066
rect 5176 19014 5228 19066
rect 5240 19014 5292 19066
rect 5304 19014 5356 19066
rect 5368 19014 5420 19066
rect 9827 19014 9879 19066
rect 9891 19014 9943 19066
rect 9955 19014 10007 19066
rect 10019 19014 10071 19066
rect 10083 19014 10135 19066
rect 14542 19014 14594 19066
rect 14606 19014 14658 19066
rect 14670 19014 14722 19066
rect 14734 19014 14786 19066
rect 14798 19014 14850 19066
rect 19257 19014 19309 19066
rect 19321 19014 19373 19066
rect 19385 19014 19437 19066
rect 19449 19014 19501 19066
rect 19513 19014 19565 19066
rect 17408 18912 17460 18964
rect 16580 18751 16632 18760
rect 16580 18717 16589 18751
rect 16589 18717 16623 18751
rect 16623 18717 16632 18751
rect 16580 18708 16632 18717
rect 18328 18751 18380 18760
rect 18328 18717 18337 18751
rect 18337 18717 18371 18751
rect 18371 18717 18380 18751
rect 18328 18708 18380 18717
rect 17316 18615 17368 18624
rect 17316 18581 17325 18615
rect 17325 18581 17359 18615
rect 17359 18581 17368 18615
rect 17316 18572 17368 18581
rect 17684 18615 17736 18624
rect 17684 18581 17693 18615
rect 17693 18581 17727 18615
rect 17727 18581 17736 18615
rect 17684 18572 17736 18581
rect 2755 18470 2807 18522
rect 2819 18470 2871 18522
rect 2883 18470 2935 18522
rect 2947 18470 2999 18522
rect 3011 18470 3063 18522
rect 7470 18470 7522 18522
rect 7534 18470 7586 18522
rect 7598 18470 7650 18522
rect 7662 18470 7714 18522
rect 7726 18470 7778 18522
rect 12185 18470 12237 18522
rect 12249 18470 12301 18522
rect 12313 18470 12365 18522
rect 12377 18470 12429 18522
rect 12441 18470 12493 18522
rect 16900 18470 16952 18522
rect 16964 18470 17016 18522
rect 17028 18470 17080 18522
rect 17092 18470 17144 18522
rect 17156 18470 17208 18522
rect 17684 18368 17736 18420
rect 18328 18368 18380 18420
rect 16580 18275 16632 18284
rect 16580 18241 16589 18275
rect 16589 18241 16623 18275
rect 16623 18241 16632 18275
rect 16580 18232 16632 18241
rect 14096 18164 14148 18216
rect 5112 17926 5164 17978
rect 5176 17926 5228 17978
rect 5240 17926 5292 17978
rect 5304 17926 5356 17978
rect 5368 17926 5420 17978
rect 9827 17926 9879 17978
rect 9891 17926 9943 17978
rect 9955 17926 10007 17978
rect 10019 17926 10071 17978
rect 10083 17926 10135 17978
rect 14542 17926 14594 17978
rect 14606 17926 14658 17978
rect 14670 17926 14722 17978
rect 14734 17926 14786 17978
rect 14798 17926 14850 17978
rect 19257 17926 19309 17978
rect 19321 17926 19373 17978
rect 19385 17926 19437 17978
rect 19449 17926 19501 17978
rect 19513 17926 19565 17978
rect 19064 17799 19116 17808
rect 19064 17765 19073 17799
rect 19073 17765 19107 17799
rect 19107 17765 19116 17799
rect 19064 17756 19116 17765
rect 17592 17527 17644 17536
rect 17592 17493 17601 17527
rect 17601 17493 17635 17527
rect 17635 17493 17644 17527
rect 17592 17484 17644 17493
rect 2755 17382 2807 17434
rect 2819 17382 2871 17434
rect 2883 17382 2935 17434
rect 2947 17382 2999 17434
rect 3011 17382 3063 17434
rect 7470 17382 7522 17434
rect 7534 17382 7586 17434
rect 7598 17382 7650 17434
rect 7662 17382 7714 17434
rect 7726 17382 7778 17434
rect 12185 17382 12237 17434
rect 12249 17382 12301 17434
rect 12313 17382 12365 17434
rect 12377 17382 12429 17434
rect 12441 17382 12493 17434
rect 16900 17382 16952 17434
rect 16964 17382 17016 17434
rect 17028 17382 17080 17434
rect 17092 17382 17144 17434
rect 17156 17382 17208 17434
rect 1216 17212 1268 17264
rect 17316 17144 17368 17196
rect 18604 17076 18656 17128
rect 5112 16838 5164 16890
rect 5176 16838 5228 16890
rect 5240 16838 5292 16890
rect 5304 16838 5356 16890
rect 5368 16838 5420 16890
rect 9827 16838 9879 16890
rect 9891 16838 9943 16890
rect 9955 16838 10007 16890
rect 10019 16838 10071 16890
rect 10083 16838 10135 16890
rect 14542 16838 14594 16890
rect 14606 16838 14658 16890
rect 14670 16838 14722 16890
rect 14734 16838 14786 16890
rect 14798 16838 14850 16890
rect 19257 16838 19309 16890
rect 19321 16838 19373 16890
rect 19385 16838 19437 16890
rect 19449 16838 19501 16890
rect 19513 16838 19565 16890
rect 14096 16779 14148 16788
rect 14096 16745 14105 16779
rect 14105 16745 14139 16779
rect 14139 16745 14148 16779
rect 14096 16736 14148 16745
rect 17592 16736 17644 16788
rect 18604 16779 18656 16788
rect 18604 16745 18613 16779
rect 18613 16745 18647 16779
rect 18647 16745 18656 16779
rect 18604 16736 18656 16745
rect 2755 16294 2807 16346
rect 2819 16294 2871 16346
rect 2883 16294 2935 16346
rect 2947 16294 2999 16346
rect 3011 16294 3063 16346
rect 7470 16294 7522 16346
rect 7534 16294 7586 16346
rect 7598 16294 7650 16346
rect 7662 16294 7714 16346
rect 7726 16294 7778 16346
rect 12185 16294 12237 16346
rect 12249 16294 12301 16346
rect 12313 16294 12365 16346
rect 12377 16294 12429 16346
rect 12441 16294 12493 16346
rect 16900 16294 16952 16346
rect 16964 16294 17016 16346
rect 17028 16294 17080 16346
rect 17092 16294 17144 16346
rect 17156 16294 17208 16346
rect 5112 15750 5164 15802
rect 5176 15750 5228 15802
rect 5240 15750 5292 15802
rect 5304 15750 5356 15802
rect 5368 15750 5420 15802
rect 9827 15750 9879 15802
rect 9891 15750 9943 15802
rect 9955 15750 10007 15802
rect 10019 15750 10071 15802
rect 10083 15750 10135 15802
rect 14542 15750 14594 15802
rect 14606 15750 14658 15802
rect 14670 15750 14722 15802
rect 14734 15750 14786 15802
rect 14798 15750 14850 15802
rect 19257 15750 19309 15802
rect 19321 15750 19373 15802
rect 19385 15750 19437 15802
rect 19449 15750 19501 15802
rect 19513 15750 19565 15802
rect 2755 15206 2807 15258
rect 2819 15206 2871 15258
rect 2883 15206 2935 15258
rect 2947 15206 2999 15258
rect 3011 15206 3063 15258
rect 7470 15206 7522 15258
rect 7534 15206 7586 15258
rect 7598 15206 7650 15258
rect 7662 15206 7714 15258
rect 7726 15206 7778 15258
rect 12185 15206 12237 15258
rect 12249 15206 12301 15258
rect 12313 15206 12365 15258
rect 12377 15206 12429 15258
rect 12441 15206 12493 15258
rect 16900 15206 16952 15258
rect 16964 15206 17016 15258
rect 17028 15206 17080 15258
rect 17092 15206 17144 15258
rect 17156 15206 17208 15258
rect 5112 14662 5164 14714
rect 5176 14662 5228 14714
rect 5240 14662 5292 14714
rect 5304 14662 5356 14714
rect 5368 14662 5420 14714
rect 9827 14662 9879 14714
rect 9891 14662 9943 14714
rect 9955 14662 10007 14714
rect 10019 14662 10071 14714
rect 10083 14662 10135 14714
rect 14542 14662 14594 14714
rect 14606 14662 14658 14714
rect 14670 14662 14722 14714
rect 14734 14662 14786 14714
rect 14798 14662 14850 14714
rect 19257 14662 19309 14714
rect 19321 14662 19373 14714
rect 19385 14662 19437 14714
rect 19449 14662 19501 14714
rect 19513 14662 19565 14714
rect 2755 14118 2807 14170
rect 2819 14118 2871 14170
rect 2883 14118 2935 14170
rect 2947 14118 2999 14170
rect 3011 14118 3063 14170
rect 7470 14118 7522 14170
rect 7534 14118 7586 14170
rect 7598 14118 7650 14170
rect 7662 14118 7714 14170
rect 7726 14118 7778 14170
rect 12185 14118 12237 14170
rect 12249 14118 12301 14170
rect 12313 14118 12365 14170
rect 12377 14118 12429 14170
rect 12441 14118 12493 14170
rect 16900 14118 16952 14170
rect 16964 14118 17016 14170
rect 17028 14118 17080 14170
rect 17092 14118 17144 14170
rect 17156 14118 17208 14170
rect 5112 13574 5164 13626
rect 5176 13574 5228 13626
rect 5240 13574 5292 13626
rect 5304 13574 5356 13626
rect 5368 13574 5420 13626
rect 9827 13574 9879 13626
rect 9891 13574 9943 13626
rect 9955 13574 10007 13626
rect 10019 13574 10071 13626
rect 10083 13574 10135 13626
rect 14542 13574 14594 13626
rect 14606 13574 14658 13626
rect 14670 13574 14722 13626
rect 14734 13574 14786 13626
rect 14798 13574 14850 13626
rect 19257 13574 19309 13626
rect 19321 13574 19373 13626
rect 19385 13574 19437 13626
rect 19449 13574 19501 13626
rect 19513 13574 19565 13626
rect 2755 13030 2807 13082
rect 2819 13030 2871 13082
rect 2883 13030 2935 13082
rect 2947 13030 2999 13082
rect 3011 13030 3063 13082
rect 7470 13030 7522 13082
rect 7534 13030 7586 13082
rect 7598 13030 7650 13082
rect 7662 13030 7714 13082
rect 7726 13030 7778 13082
rect 12185 13030 12237 13082
rect 12249 13030 12301 13082
rect 12313 13030 12365 13082
rect 12377 13030 12429 13082
rect 12441 13030 12493 13082
rect 16900 13030 16952 13082
rect 16964 13030 17016 13082
rect 17028 13030 17080 13082
rect 17092 13030 17144 13082
rect 17156 13030 17208 13082
rect 5112 12486 5164 12538
rect 5176 12486 5228 12538
rect 5240 12486 5292 12538
rect 5304 12486 5356 12538
rect 5368 12486 5420 12538
rect 9827 12486 9879 12538
rect 9891 12486 9943 12538
rect 9955 12486 10007 12538
rect 10019 12486 10071 12538
rect 10083 12486 10135 12538
rect 14542 12486 14594 12538
rect 14606 12486 14658 12538
rect 14670 12486 14722 12538
rect 14734 12486 14786 12538
rect 14798 12486 14850 12538
rect 19257 12486 19309 12538
rect 19321 12486 19373 12538
rect 19385 12486 19437 12538
rect 19449 12486 19501 12538
rect 19513 12486 19565 12538
rect 2755 11942 2807 11994
rect 2819 11942 2871 11994
rect 2883 11942 2935 11994
rect 2947 11942 2999 11994
rect 3011 11942 3063 11994
rect 7470 11942 7522 11994
rect 7534 11942 7586 11994
rect 7598 11942 7650 11994
rect 7662 11942 7714 11994
rect 7726 11942 7778 11994
rect 12185 11942 12237 11994
rect 12249 11942 12301 11994
rect 12313 11942 12365 11994
rect 12377 11942 12429 11994
rect 12441 11942 12493 11994
rect 16900 11942 16952 11994
rect 16964 11942 17016 11994
rect 17028 11942 17080 11994
rect 17092 11942 17144 11994
rect 17156 11942 17208 11994
rect 5112 11398 5164 11450
rect 5176 11398 5228 11450
rect 5240 11398 5292 11450
rect 5304 11398 5356 11450
rect 5368 11398 5420 11450
rect 9827 11398 9879 11450
rect 9891 11398 9943 11450
rect 9955 11398 10007 11450
rect 10019 11398 10071 11450
rect 10083 11398 10135 11450
rect 14542 11398 14594 11450
rect 14606 11398 14658 11450
rect 14670 11398 14722 11450
rect 14734 11398 14786 11450
rect 14798 11398 14850 11450
rect 19257 11398 19309 11450
rect 19321 11398 19373 11450
rect 19385 11398 19437 11450
rect 19449 11398 19501 11450
rect 19513 11398 19565 11450
rect 2755 10854 2807 10906
rect 2819 10854 2871 10906
rect 2883 10854 2935 10906
rect 2947 10854 2999 10906
rect 3011 10854 3063 10906
rect 7470 10854 7522 10906
rect 7534 10854 7586 10906
rect 7598 10854 7650 10906
rect 7662 10854 7714 10906
rect 7726 10854 7778 10906
rect 12185 10854 12237 10906
rect 12249 10854 12301 10906
rect 12313 10854 12365 10906
rect 12377 10854 12429 10906
rect 12441 10854 12493 10906
rect 16900 10854 16952 10906
rect 16964 10854 17016 10906
rect 17028 10854 17080 10906
rect 17092 10854 17144 10906
rect 17156 10854 17208 10906
rect 5112 10310 5164 10362
rect 5176 10310 5228 10362
rect 5240 10310 5292 10362
rect 5304 10310 5356 10362
rect 5368 10310 5420 10362
rect 9827 10310 9879 10362
rect 9891 10310 9943 10362
rect 9955 10310 10007 10362
rect 10019 10310 10071 10362
rect 10083 10310 10135 10362
rect 14542 10310 14594 10362
rect 14606 10310 14658 10362
rect 14670 10310 14722 10362
rect 14734 10310 14786 10362
rect 14798 10310 14850 10362
rect 19257 10310 19309 10362
rect 19321 10310 19373 10362
rect 19385 10310 19437 10362
rect 19449 10310 19501 10362
rect 19513 10310 19565 10362
rect 19064 9911 19116 9920
rect 19064 9877 19073 9911
rect 19073 9877 19107 9911
rect 19107 9877 19116 9911
rect 19064 9868 19116 9877
rect 2755 9766 2807 9818
rect 2819 9766 2871 9818
rect 2883 9766 2935 9818
rect 2947 9766 2999 9818
rect 3011 9766 3063 9818
rect 7470 9766 7522 9818
rect 7534 9766 7586 9818
rect 7598 9766 7650 9818
rect 7662 9766 7714 9818
rect 7726 9766 7778 9818
rect 12185 9766 12237 9818
rect 12249 9766 12301 9818
rect 12313 9766 12365 9818
rect 12377 9766 12429 9818
rect 12441 9766 12493 9818
rect 16900 9766 16952 9818
rect 16964 9766 17016 9818
rect 17028 9766 17080 9818
rect 17092 9766 17144 9818
rect 17156 9766 17208 9818
rect 5112 9222 5164 9274
rect 5176 9222 5228 9274
rect 5240 9222 5292 9274
rect 5304 9222 5356 9274
rect 5368 9222 5420 9274
rect 9827 9222 9879 9274
rect 9891 9222 9943 9274
rect 9955 9222 10007 9274
rect 10019 9222 10071 9274
rect 10083 9222 10135 9274
rect 14542 9222 14594 9274
rect 14606 9222 14658 9274
rect 14670 9222 14722 9274
rect 14734 9222 14786 9274
rect 14798 9222 14850 9274
rect 19257 9222 19309 9274
rect 19321 9222 19373 9274
rect 19385 9222 19437 9274
rect 19449 9222 19501 9274
rect 19513 9222 19565 9274
rect 2755 8678 2807 8730
rect 2819 8678 2871 8730
rect 2883 8678 2935 8730
rect 2947 8678 2999 8730
rect 3011 8678 3063 8730
rect 7470 8678 7522 8730
rect 7534 8678 7586 8730
rect 7598 8678 7650 8730
rect 7662 8678 7714 8730
rect 7726 8678 7778 8730
rect 12185 8678 12237 8730
rect 12249 8678 12301 8730
rect 12313 8678 12365 8730
rect 12377 8678 12429 8730
rect 12441 8678 12493 8730
rect 16900 8678 16952 8730
rect 16964 8678 17016 8730
rect 17028 8678 17080 8730
rect 17092 8678 17144 8730
rect 17156 8678 17208 8730
rect 5112 8134 5164 8186
rect 5176 8134 5228 8186
rect 5240 8134 5292 8186
rect 5304 8134 5356 8186
rect 5368 8134 5420 8186
rect 9827 8134 9879 8186
rect 9891 8134 9943 8186
rect 9955 8134 10007 8186
rect 10019 8134 10071 8186
rect 10083 8134 10135 8186
rect 14542 8134 14594 8186
rect 14606 8134 14658 8186
rect 14670 8134 14722 8186
rect 14734 8134 14786 8186
rect 14798 8134 14850 8186
rect 19257 8134 19309 8186
rect 19321 8134 19373 8186
rect 19385 8134 19437 8186
rect 19449 8134 19501 8186
rect 19513 8134 19565 8186
rect 2755 7590 2807 7642
rect 2819 7590 2871 7642
rect 2883 7590 2935 7642
rect 2947 7590 2999 7642
rect 3011 7590 3063 7642
rect 7470 7590 7522 7642
rect 7534 7590 7586 7642
rect 7598 7590 7650 7642
rect 7662 7590 7714 7642
rect 7726 7590 7778 7642
rect 12185 7590 12237 7642
rect 12249 7590 12301 7642
rect 12313 7590 12365 7642
rect 12377 7590 12429 7642
rect 12441 7590 12493 7642
rect 16900 7590 16952 7642
rect 16964 7590 17016 7642
rect 17028 7590 17080 7642
rect 17092 7590 17144 7642
rect 17156 7590 17208 7642
rect 5112 7046 5164 7098
rect 5176 7046 5228 7098
rect 5240 7046 5292 7098
rect 5304 7046 5356 7098
rect 5368 7046 5420 7098
rect 9827 7046 9879 7098
rect 9891 7046 9943 7098
rect 9955 7046 10007 7098
rect 10019 7046 10071 7098
rect 10083 7046 10135 7098
rect 14542 7046 14594 7098
rect 14606 7046 14658 7098
rect 14670 7046 14722 7098
rect 14734 7046 14786 7098
rect 14798 7046 14850 7098
rect 19257 7046 19309 7098
rect 19321 7046 19373 7098
rect 19385 7046 19437 7098
rect 19449 7046 19501 7098
rect 19513 7046 19565 7098
rect 2755 6502 2807 6554
rect 2819 6502 2871 6554
rect 2883 6502 2935 6554
rect 2947 6502 2999 6554
rect 3011 6502 3063 6554
rect 7470 6502 7522 6554
rect 7534 6502 7586 6554
rect 7598 6502 7650 6554
rect 7662 6502 7714 6554
rect 7726 6502 7778 6554
rect 12185 6502 12237 6554
rect 12249 6502 12301 6554
rect 12313 6502 12365 6554
rect 12377 6502 12429 6554
rect 12441 6502 12493 6554
rect 16900 6502 16952 6554
rect 16964 6502 17016 6554
rect 17028 6502 17080 6554
rect 17092 6502 17144 6554
rect 17156 6502 17208 6554
rect 5112 5958 5164 6010
rect 5176 5958 5228 6010
rect 5240 5958 5292 6010
rect 5304 5958 5356 6010
rect 5368 5958 5420 6010
rect 9827 5958 9879 6010
rect 9891 5958 9943 6010
rect 9955 5958 10007 6010
rect 10019 5958 10071 6010
rect 10083 5958 10135 6010
rect 14542 5958 14594 6010
rect 14606 5958 14658 6010
rect 14670 5958 14722 6010
rect 14734 5958 14786 6010
rect 14798 5958 14850 6010
rect 19257 5958 19309 6010
rect 19321 5958 19373 6010
rect 19385 5958 19437 6010
rect 19449 5958 19501 6010
rect 19513 5958 19565 6010
rect 2755 5414 2807 5466
rect 2819 5414 2871 5466
rect 2883 5414 2935 5466
rect 2947 5414 2999 5466
rect 3011 5414 3063 5466
rect 7470 5414 7522 5466
rect 7534 5414 7586 5466
rect 7598 5414 7650 5466
rect 7662 5414 7714 5466
rect 7726 5414 7778 5466
rect 12185 5414 12237 5466
rect 12249 5414 12301 5466
rect 12313 5414 12365 5466
rect 12377 5414 12429 5466
rect 12441 5414 12493 5466
rect 16900 5414 16952 5466
rect 16964 5414 17016 5466
rect 17028 5414 17080 5466
rect 17092 5414 17144 5466
rect 17156 5414 17208 5466
rect 5112 4870 5164 4922
rect 5176 4870 5228 4922
rect 5240 4870 5292 4922
rect 5304 4870 5356 4922
rect 5368 4870 5420 4922
rect 9827 4870 9879 4922
rect 9891 4870 9943 4922
rect 9955 4870 10007 4922
rect 10019 4870 10071 4922
rect 10083 4870 10135 4922
rect 14542 4870 14594 4922
rect 14606 4870 14658 4922
rect 14670 4870 14722 4922
rect 14734 4870 14786 4922
rect 14798 4870 14850 4922
rect 19257 4870 19309 4922
rect 19321 4870 19373 4922
rect 19385 4870 19437 4922
rect 19449 4870 19501 4922
rect 19513 4870 19565 4922
rect 2755 4326 2807 4378
rect 2819 4326 2871 4378
rect 2883 4326 2935 4378
rect 2947 4326 2999 4378
rect 3011 4326 3063 4378
rect 7470 4326 7522 4378
rect 7534 4326 7586 4378
rect 7598 4326 7650 4378
rect 7662 4326 7714 4378
rect 7726 4326 7778 4378
rect 12185 4326 12237 4378
rect 12249 4326 12301 4378
rect 12313 4326 12365 4378
rect 12377 4326 12429 4378
rect 12441 4326 12493 4378
rect 16900 4326 16952 4378
rect 16964 4326 17016 4378
rect 17028 4326 17080 4378
rect 17092 4326 17144 4378
rect 17156 4326 17208 4378
rect 5112 3782 5164 3834
rect 5176 3782 5228 3834
rect 5240 3782 5292 3834
rect 5304 3782 5356 3834
rect 5368 3782 5420 3834
rect 9827 3782 9879 3834
rect 9891 3782 9943 3834
rect 9955 3782 10007 3834
rect 10019 3782 10071 3834
rect 10083 3782 10135 3834
rect 14542 3782 14594 3834
rect 14606 3782 14658 3834
rect 14670 3782 14722 3834
rect 14734 3782 14786 3834
rect 14798 3782 14850 3834
rect 19257 3782 19309 3834
rect 19321 3782 19373 3834
rect 19385 3782 19437 3834
rect 19449 3782 19501 3834
rect 19513 3782 19565 3834
rect 2755 3238 2807 3290
rect 2819 3238 2871 3290
rect 2883 3238 2935 3290
rect 2947 3238 2999 3290
rect 3011 3238 3063 3290
rect 7470 3238 7522 3290
rect 7534 3238 7586 3290
rect 7598 3238 7650 3290
rect 7662 3238 7714 3290
rect 7726 3238 7778 3290
rect 12185 3238 12237 3290
rect 12249 3238 12301 3290
rect 12313 3238 12365 3290
rect 12377 3238 12429 3290
rect 12441 3238 12493 3290
rect 16900 3238 16952 3290
rect 16964 3238 17016 3290
rect 17028 3238 17080 3290
rect 17092 3238 17144 3290
rect 17156 3238 17208 3290
rect 5112 2694 5164 2746
rect 5176 2694 5228 2746
rect 5240 2694 5292 2746
rect 5304 2694 5356 2746
rect 5368 2694 5420 2746
rect 9827 2694 9879 2746
rect 9891 2694 9943 2746
rect 9955 2694 10007 2746
rect 10019 2694 10071 2746
rect 10083 2694 10135 2746
rect 14542 2694 14594 2746
rect 14606 2694 14658 2746
rect 14670 2694 14722 2746
rect 14734 2694 14786 2746
rect 14798 2694 14850 2746
rect 19257 2694 19309 2746
rect 19321 2694 19373 2746
rect 19385 2694 19437 2746
rect 19449 2694 19501 2746
rect 19513 2694 19565 2746
rect 2755 2150 2807 2202
rect 2819 2150 2871 2202
rect 2883 2150 2935 2202
rect 2947 2150 2999 2202
rect 3011 2150 3063 2202
rect 7470 2150 7522 2202
rect 7534 2150 7586 2202
rect 7598 2150 7650 2202
rect 7662 2150 7714 2202
rect 7726 2150 7778 2202
rect 12185 2150 12237 2202
rect 12249 2150 12301 2202
rect 12313 2150 12365 2202
rect 12377 2150 12429 2202
rect 12441 2150 12493 2202
rect 16900 2150 16952 2202
rect 16964 2150 17016 2202
rect 17028 2150 17080 2202
rect 17092 2150 17144 2202
rect 17156 2150 17208 2202
rect 5112 1606 5164 1658
rect 5176 1606 5228 1658
rect 5240 1606 5292 1658
rect 5304 1606 5356 1658
rect 5368 1606 5420 1658
rect 9827 1606 9879 1658
rect 9891 1606 9943 1658
rect 9955 1606 10007 1658
rect 10019 1606 10071 1658
rect 10083 1606 10135 1658
rect 14542 1606 14594 1658
rect 14606 1606 14658 1658
rect 14670 1606 14722 1658
rect 14734 1606 14786 1658
rect 14798 1606 14850 1658
rect 19257 1606 19309 1658
rect 19321 1606 19373 1658
rect 19385 1606 19437 1658
rect 19449 1606 19501 1658
rect 19513 1606 19565 1658
rect 2755 1062 2807 1114
rect 2819 1062 2871 1114
rect 2883 1062 2935 1114
rect 2947 1062 2999 1114
rect 3011 1062 3063 1114
rect 7470 1062 7522 1114
rect 7534 1062 7586 1114
rect 7598 1062 7650 1114
rect 7662 1062 7714 1114
rect 7726 1062 7778 1114
rect 12185 1062 12237 1114
rect 12249 1062 12301 1114
rect 12313 1062 12365 1114
rect 12377 1062 12429 1114
rect 12441 1062 12493 1114
rect 16900 1062 16952 1114
rect 16964 1062 17016 1114
rect 17028 1062 17080 1114
rect 17092 1062 17144 1114
rect 17156 1062 17208 1114
rect 3792 799 3844 808
rect 3792 765 3801 799
rect 3801 765 3835 799
rect 3835 765 3844 799
rect 3792 756 3844 765
rect 6276 799 6328 808
rect 6276 765 6285 799
rect 6285 765 6319 799
rect 6319 765 6328 799
rect 6276 756 6328 765
rect 8760 799 8812 808
rect 8760 765 8769 799
rect 8769 765 8803 799
rect 8803 765 8812 799
rect 8760 756 8812 765
rect 11244 799 11296 808
rect 11244 765 11253 799
rect 11253 765 11287 799
rect 11287 765 11296 799
rect 11244 756 11296 765
rect 13728 799 13780 808
rect 13728 765 13737 799
rect 13737 765 13771 799
rect 13771 765 13780 799
rect 13728 756 13780 765
rect 16212 799 16264 808
rect 16212 765 16221 799
rect 16221 765 16255 799
rect 16255 765 16264 799
rect 16212 756 16264 765
rect 18696 799 18748 808
rect 18696 765 18705 799
rect 18705 765 18739 799
rect 18739 765 18748 799
rect 18696 756 18748 765
rect 5112 518 5164 570
rect 5176 518 5228 570
rect 5240 518 5292 570
rect 5304 518 5356 570
rect 5368 518 5420 570
rect 9827 518 9879 570
rect 9891 518 9943 570
rect 9955 518 10007 570
rect 10019 518 10071 570
rect 10083 518 10135 570
rect 14542 518 14594 570
rect 14606 518 14658 570
rect 14670 518 14722 570
rect 14734 518 14786 570
rect 14798 518 14850 570
rect 19257 518 19309 570
rect 19321 518 19373 570
rect 19385 518 19437 570
rect 19449 518 19501 570
rect 19513 518 19565 570
<< metal2 >>
rect 846 19600 902 20000
rect 2502 19600 2558 20000
rect 4158 19600 4214 20000
rect 5814 19600 5870 20000
rect 7470 19600 7526 20000
rect 9126 19600 9182 20000
rect 10782 19600 10838 20000
rect 12438 19600 12494 20000
rect 14094 19600 14150 20000
rect 15750 19600 15806 20000
rect 17406 19600 17462 20000
rect 19062 19600 19118 20000
rect 5112 19068 5420 19077
rect 5112 19066 5118 19068
rect 5174 19066 5198 19068
rect 5254 19066 5278 19068
rect 5334 19066 5358 19068
rect 5414 19066 5420 19068
rect 5174 19014 5176 19066
rect 5356 19014 5358 19066
rect 5112 19012 5118 19014
rect 5174 19012 5198 19014
rect 5254 19012 5278 19014
rect 5334 19012 5358 19014
rect 5414 19012 5420 19014
rect 5112 19003 5420 19012
rect 9827 19068 10135 19077
rect 9827 19066 9833 19068
rect 9889 19066 9913 19068
rect 9969 19066 9993 19068
rect 10049 19066 10073 19068
rect 10129 19066 10135 19068
rect 9889 19014 9891 19066
rect 10071 19014 10073 19066
rect 9827 19012 9833 19014
rect 9889 19012 9913 19014
rect 9969 19012 9993 19014
rect 10049 19012 10073 19014
rect 10129 19012 10135 19014
rect 9827 19003 10135 19012
rect 14542 19068 14850 19077
rect 14542 19066 14548 19068
rect 14604 19066 14628 19068
rect 14684 19066 14708 19068
rect 14764 19066 14788 19068
rect 14844 19066 14850 19068
rect 14604 19014 14606 19066
rect 14786 19014 14788 19066
rect 14542 19012 14548 19014
rect 14604 19012 14628 19014
rect 14684 19012 14708 19014
rect 14764 19012 14788 19014
rect 14844 19012 14850 19014
rect 14542 19003 14850 19012
rect 17420 18970 17448 19600
rect 17408 18964 17460 18970
rect 17408 18906 17460 18912
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 2755 18524 3063 18533
rect 2755 18522 2761 18524
rect 2817 18522 2841 18524
rect 2897 18522 2921 18524
rect 2977 18522 3001 18524
rect 3057 18522 3063 18524
rect 2817 18470 2819 18522
rect 2999 18470 3001 18522
rect 2755 18468 2761 18470
rect 2817 18468 2841 18470
rect 2897 18468 2921 18470
rect 2977 18468 3001 18470
rect 3057 18468 3063 18470
rect 2755 18459 3063 18468
rect 7470 18524 7778 18533
rect 7470 18522 7476 18524
rect 7532 18522 7556 18524
rect 7612 18522 7636 18524
rect 7692 18522 7716 18524
rect 7772 18522 7778 18524
rect 7532 18470 7534 18522
rect 7714 18470 7716 18522
rect 7470 18468 7476 18470
rect 7532 18468 7556 18470
rect 7612 18468 7636 18470
rect 7692 18468 7716 18470
rect 7772 18468 7778 18470
rect 7470 18459 7778 18468
rect 12185 18524 12493 18533
rect 12185 18522 12191 18524
rect 12247 18522 12271 18524
rect 12327 18522 12351 18524
rect 12407 18522 12431 18524
rect 12487 18522 12493 18524
rect 12247 18470 12249 18522
rect 12429 18470 12431 18522
rect 12185 18468 12191 18470
rect 12247 18468 12271 18470
rect 12327 18468 12351 18470
rect 12407 18468 12431 18470
rect 12487 18468 12493 18470
rect 12185 18459 12493 18468
rect 16592 18290 16620 18702
rect 17316 18624 17368 18630
rect 17316 18566 17368 18572
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 16900 18524 17208 18533
rect 16900 18522 16906 18524
rect 16962 18522 16986 18524
rect 17042 18522 17066 18524
rect 17122 18522 17146 18524
rect 17202 18522 17208 18524
rect 16962 18470 16964 18522
rect 17144 18470 17146 18522
rect 16900 18468 16906 18470
rect 16962 18468 16986 18470
rect 17042 18468 17066 18470
rect 17122 18468 17146 18470
rect 17202 18468 17208 18470
rect 16900 18459 17208 18468
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 5112 17980 5420 17989
rect 5112 17978 5118 17980
rect 5174 17978 5198 17980
rect 5254 17978 5278 17980
rect 5334 17978 5358 17980
rect 5414 17978 5420 17980
rect 5174 17926 5176 17978
rect 5356 17926 5358 17978
rect 5112 17924 5118 17926
rect 5174 17924 5198 17926
rect 5254 17924 5278 17926
rect 5334 17924 5358 17926
rect 5414 17924 5420 17926
rect 5112 17915 5420 17924
rect 9827 17980 10135 17989
rect 9827 17978 9833 17980
rect 9889 17978 9913 17980
rect 9969 17978 9993 17980
rect 10049 17978 10073 17980
rect 10129 17978 10135 17980
rect 9889 17926 9891 17978
rect 10071 17926 10073 17978
rect 9827 17924 9833 17926
rect 9889 17924 9913 17926
rect 9969 17924 9993 17926
rect 10049 17924 10073 17926
rect 10129 17924 10135 17926
rect 9827 17915 10135 17924
rect 2755 17436 3063 17445
rect 2755 17434 2761 17436
rect 2817 17434 2841 17436
rect 2897 17434 2921 17436
rect 2977 17434 3001 17436
rect 3057 17434 3063 17436
rect 2817 17382 2819 17434
rect 2999 17382 3001 17434
rect 2755 17380 2761 17382
rect 2817 17380 2841 17382
rect 2897 17380 2921 17382
rect 2977 17380 3001 17382
rect 3057 17380 3063 17382
rect 2755 17371 3063 17380
rect 7470 17436 7778 17445
rect 7470 17434 7476 17436
rect 7532 17434 7556 17436
rect 7612 17434 7636 17436
rect 7692 17434 7716 17436
rect 7772 17434 7778 17436
rect 7532 17382 7534 17434
rect 7714 17382 7716 17434
rect 7470 17380 7476 17382
rect 7532 17380 7556 17382
rect 7612 17380 7636 17382
rect 7692 17380 7716 17382
rect 7772 17380 7778 17382
rect 7470 17371 7778 17380
rect 12185 17436 12493 17445
rect 12185 17434 12191 17436
rect 12247 17434 12271 17436
rect 12327 17434 12351 17436
rect 12407 17434 12431 17436
rect 12487 17434 12493 17436
rect 12247 17382 12249 17434
rect 12429 17382 12431 17434
rect 12185 17380 12191 17382
rect 12247 17380 12271 17382
rect 12327 17380 12351 17382
rect 12407 17380 12431 17382
rect 12487 17380 12493 17382
rect 12185 17371 12493 17380
rect 1216 17264 1268 17270
rect 1216 17206 1268 17212
rect 1228 400 1256 17206
rect 5112 16892 5420 16901
rect 5112 16890 5118 16892
rect 5174 16890 5198 16892
rect 5254 16890 5278 16892
rect 5334 16890 5358 16892
rect 5414 16890 5420 16892
rect 5174 16838 5176 16890
rect 5356 16838 5358 16890
rect 5112 16836 5118 16838
rect 5174 16836 5198 16838
rect 5254 16836 5278 16838
rect 5334 16836 5358 16838
rect 5414 16836 5420 16838
rect 5112 16827 5420 16836
rect 9827 16892 10135 16901
rect 9827 16890 9833 16892
rect 9889 16890 9913 16892
rect 9969 16890 9993 16892
rect 10049 16890 10073 16892
rect 10129 16890 10135 16892
rect 9889 16838 9891 16890
rect 10071 16838 10073 16890
rect 9827 16836 9833 16838
rect 9889 16836 9913 16838
rect 9969 16836 9993 16838
rect 10049 16836 10073 16838
rect 10129 16836 10135 16838
rect 9827 16827 10135 16836
rect 14108 16794 14136 18158
rect 14542 17980 14850 17989
rect 14542 17978 14548 17980
rect 14604 17978 14628 17980
rect 14684 17978 14708 17980
rect 14764 17978 14788 17980
rect 14844 17978 14850 17980
rect 14604 17926 14606 17978
rect 14786 17926 14788 17978
rect 14542 17924 14548 17926
rect 14604 17924 14628 17926
rect 14684 17924 14708 17926
rect 14764 17924 14788 17926
rect 14844 17924 14850 17926
rect 14542 17915 14850 17924
rect 16900 17436 17208 17445
rect 16900 17434 16906 17436
rect 16962 17434 16986 17436
rect 17042 17434 17066 17436
rect 17122 17434 17146 17436
rect 17202 17434 17208 17436
rect 16962 17382 16964 17434
rect 17144 17382 17146 17434
rect 16900 17380 16906 17382
rect 16962 17380 16986 17382
rect 17042 17380 17066 17382
rect 17122 17380 17146 17382
rect 17202 17380 17208 17382
rect 16900 17371 17208 17380
rect 17328 17202 17356 18566
rect 17696 18426 17724 18566
rect 18340 18426 18368 18702
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 19076 17814 19104 19600
rect 19257 19068 19565 19077
rect 19257 19066 19263 19068
rect 19319 19066 19343 19068
rect 19399 19066 19423 19068
rect 19479 19066 19503 19068
rect 19559 19066 19565 19068
rect 19319 19014 19321 19066
rect 19501 19014 19503 19066
rect 19257 19012 19263 19014
rect 19319 19012 19343 19014
rect 19399 19012 19423 19014
rect 19479 19012 19503 19014
rect 19559 19012 19565 19014
rect 19257 19003 19565 19012
rect 19257 17980 19565 17989
rect 19257 17978 19263 17980
rect 19319 17978 19343 17980
rect 19399 17978 19423 17980
rect 19479 17978 19503 17980
rect 19559 17978 19565 17980
rect 19319 17926 19321 17978
rect 19501 17926 19503 17978
rect 19257 17924 19263 17926
rect 19319 17924 19343 17926
rect 19399 17924 19423 17926
rect 19479 17924 19503 17926
rect 19559 17924 19565 17926
rect 19257 17915 19565 17924
rect 19064 17808 19116 17814
rect 19064 17750 19116 17756
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 14542 16892 14850 16901
rect 14542 16890 14548 16892
rect 14604 16890 14628 16892
rect 14684 16890 14708 16892
rect 14764 16890 14788 16892
rect 14844 16890 14850 16892
rect 14604 16838 14606 16890
rect 14786 16838 14788 16890
rect 14542 16836 14548 16838
rect 14604 16836 14628 16838
rect 14684 16836 14708 16838
rect 14764 16836 14788 16838
rect 14844 16836 14850 16838
rect 14542 16827 14850 16836
rect 17604 16794 17632 17478
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18616 16794 18644 17070
rect 19257 16892 19565 16901
rect 19257 16890 19263 16892
rect 19319 16890 19343 16892
rect 19399 16890 19423 16892
rect 19479 16890 19503 16892
rect 19559 16890 19565 16892
rect 19319 16838 19321 16890
rect 19501 16838 19503 16890
rect 19257 16836 19263 16838
rect 19319 16836 19343 16838
rect 19399 16836 19423 16838
rect 19479 16836 19503 16838
rect 19559 16836 19565 16838
rect 19257 16827 19565 16836
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 2755 16348 3063 16357
rect 2755 16346 2761 16348
rect 2817 16346 2841 16348
rect 2897 16346 2921 16348
rect 2977 16346 3001 16348
rect 3057 16346 3063 16348
rect 2817 16294 2819 16346
rect 2999 16294 3001 16346
rect 2755 16292 2761 16294
rect 2817 16292 2841 16294
rect 2897 16292 2921 16294
rect 2977 16292 3001 16294
rect 3057 16292 3063 16294
rect 2755 16283 3063 16292
rect 7470 16348 7778 16357
rect 7470 16346 7476 16348
rect 7532 16346 7556 16348
rect 7612 16346 7636 16348
rect 7692 16346 7716 16348
rect 7772 16346 7778 16348
rect 7532 16294 7534 16346
rect 7714 16294 7716 16346
rect 7470 16292 7476 16294
rect 7532 16292 7556 16294
rect 7612 16292 7636 16294
rect 7692 16292 7716 16294
rect 7772 16292 7778 16294
rect 7470 16283 7778 16292
rect 12185 16348 12493 16357
rect 12185 16346 12191 16348
rect 12247 16346 12271 16348
rect 12327 16346 12351 16348
rect 12407 16346 12431 16348
rect 12487 16346 12493 16348
rect 12247 16294 12249 16346
rect 12429 16294 12431 16346
rect 12185 16292 12191 16294
rect 12247 16292 12271 16294
rect 12327 16292 12351 16294
rect 12407 16292 12431 16294
rect 12487 16292 12493 16294
rect 12185 16283 12493 16292
rect 16900 16348 17208 16357
rect 16900 16346 16906 16348
rect 16962 16346 16986 16348
rect 17042 16346 17066 16348
rect 17122 16346 17146 16348
rect 17202 16346 17208 16348
rect 16962 16294 16964 16346
rect 17144 16294 17146 16346
rect 16900 16292 16906 16294
rect 16962 16292 16986 16294
rect 17042 16292 17066 16294
rect 17122 16292 17146 16294
rect 17202 16292 17208 16294
rect 16900 16283 17208 16292
rect 5112 15804 5420 15813
rect 5112 15802 5118 15804
rect 5174 15802 5198 15804
rect 5254 15802 5278 15804
rect 5334 15802 5358 15804
rect 5414 15802 5420 15804
rect 5174 15750 5176 15802
rect 5356 15750 5358 15802
rect 5112 15748 5118 15750
rect 5174 15748 5198 15750
rect 5254 15748 5278 15750
rect 5334 15748 5358 15750
rect 5414 15748 5420 15750
rect 5112 15739 5420 15748
rect 9827 15804 10135 15813
rect 9827 15802 9833 15804
rect 9889 15802 9913 15804
rect 9969 15802 9993 15804
rect 10049 15802 10073 15804
rect 10129 15802 10135 15804
rect 9889 15750 9891 15802
rect 10071 15750 10073 15802
rect 9827 15748 9833 15750
rect 9889 15748 9913 15750
rect 9969 15748 9993 15750
rect 10049 15748 10073 15750
rect 10129 15748 10135 15750
rect 9827 15739 10135 15748
rect 14542 15804 14850 15813
rect 14542 15802 14548 15804
rect 14604 15802 14628 15804
rect 14684 15802 14708 15804
rect 14764 15802 14788 15804
rect 14844 15802 14850 15804
rect 14604 15750 14606 15802
rect 14786 15750 14788 15802
rect 14542 15748 14548 15750
rect 14604 15748 14628 15750
rect 14684 15748 14708 15750
rect 14764 15748 14788 15750
rect 14844 15748 14850 15750
rect 14542 15739 14850 15748
rect 19257 15804 19565 15813
rect 19257 15802 19263 15804
rect 19319 15802 19343 15804
rect 19399 15802 19423 15804
rect 19479 15802 19503 15804
rect 19559 15802 19565 15804
rect 19319 15750 19321 15802
rect 19501 15750 19503 15802
rect 19257 15748 19263 15750
rect 19319 15748 19343 15750
rect 19399 15748 19423 15750
rect 19479 15748 19503 15750
rect 19559 15748 19565 15750
rect 19257 15739 19565 15748
rect 2755 15260 3063 15269
rect 2755 15258 2761 15260
rect 2817 15258 2841 15260
rect 2897 15258 2921 15260
rect 2977 15258 3001 15260
rect 3057 15258 3063 15260
rect 2817 15206 2819 15258
rect 2999 15206 3001 15258
rect 2755 15204 2761 15206
rect 2817 15204 2841 15206
rect 2897 15204 2921 15206
rect 2977 15204 3001 15206
rect 3057 15204 3063 15206
rect 2755 15195 3063 15204
rect 7470 15260 7778 15269
rect 7470 15258 7476 15260
rect 7532 15258 7556 15260
rect 7612 15258 7636 15260
rect 7692 15258 7716 15260
rect 7772 15258 7778 15260
rect 7532 15206 7534 15258
rect 7714 15206 7716 15258
rect 7470 15204 7476 15206
rect 7532 15204 7556 15206
rect 7612 15204 7636 15206
rect 7692 15204 7716 15206
rect 7772 15204 7778 15206
rect 7470 15195 7778 15204
rect 12185 15260 12493 15269
rect 12185 15258 12191 15260
rect 12247 15258 12271 15260
rect 12327 15258 12351 15260
rect 12407 15258 12431 15260
rect 12487 15258 12493 15260
rect 12247 15206 12249 15258
rect 12429 15206 12431 15258
rect 12185 15204 12191 15206
rect 12247 15204 12271 15206
rect 12327 15204 12351 15206
rect 12407 15204 12431 15206
rect 12487 15204 12493 15206
rect 12185 15195 12493 15204
rect 16900 15260 17208 15269
rect 16900 15258 16906 15260
rect 16962 15258 16986 15260
rect 17042 15258 17066 15260
rect 17122 15258 17146 15260
rect 17202 15258 17208 15260
rect 16962 15206 16964 15258
rect 17144 15206 17146 15258
rect 16900 15204 16906 15206
rect 16962 15204 16986 15206
rect 17042 15204 17066 15206
rect 17122 15204 17146 15206
rect 17202 15204 17208 15206
rect 16900 15195 17208 15204
rect 5112 14716 5420 14725
rect 5112 14714 5118 14716
rect 5174 14714 5198 14716
rect 5254 14714 5278 14716
rect 5334 14714 5358 14716
rect 5414 14714 5420 14716
rect 5174 14662 5176 14714
rect 5356 14662 5358 14714
rect 5112 14660 5118 14662
rect 5174 14660 5198 14662
rect 5254 14660 5278 14662
rect 5334 14660 5358 14662
rect 5414 14660 5420 14662
rect 5112 14651 5420 14660
rect 9827 14716 10135 14725
rect 9827 14714 9833 14716
rect 9889 14714 9913 14716
rect 9969 14714 9993 14716
rect 10049 14714 10073 14716
rect 10129 14714 10135 14716
rect 9889 14662 9891 14714
rect 10071 14662 10073 14714
rect 9827 14660 9833 14662
rect 9889 14660 9913 14662
rect 9969 14660 9993 14662
rect 10049 14660 10073 14662
rect 10129 14660 10135 14662
rect 9827 14651 10135 14660
rect 14542 14716 14850 14725
rect 14542 14714 14548 14716
rect 14604 14714 14628 14716
rect 14684 14714 14708 14716
rect 14764 14714 14788 14716
rect 14844 14714 14850 14716
rect 14604 14662 14606 14714
rect 14786 14662 14788 14714
rect 14542 14660 14548 14662
rect 14604 14660 14628 14662
rect 14684 14660 14708 14662
rect 14764 14660 14788 14662
rect 14844 14660 14850 14662
rect 14542 14651 14850 14660
rect 19257 14716 19565 14725
rect 19257 14714 19263 14716
rect 19319 14714 19343 14716
rect 19399 14714 19423 14716
rect 19479 14714 19503 14716
rect 19559 14714 19565 14716
rect 19319 14662 19321 14714
rect 19501 14662 19503 14714
rect 19257 14660 19263 14662
rect 19319 14660 19343 14662
rect 19399 14660 19423 14662
rect 19479 14660 19503 14662
rect 19559 14660 19565 14662
rect 19257 14651 19565 14660
rect 2755 14172 3063 14181
rect 2755 14170 2761 14172
rect 2817 14170 2841 14172
rect 2897 14170 2921 14172
rect 2977 14170 3001 14172
rect 3057 14170 3063 14172
rect 2817 14118 2819 14170
rect 2999 14118 3001 14170
rect 2755 14116 2761 14118
rect 2817 14116 2841 14118
rect 2897 14116 2921 14118
rect 2977 14116 3001 14118
rect 3057 14116 3063 14118
rect 2755 14107 3063 14116
rect 7470 14172 7778 14181
rect 7470 14170 7476 14172
rect 7532 14170 7556 14172
rect 7612 14170 7636 14172
rect 7692 14170 7716 14172
rect 7772 14170 7778 14172
rect 7532 14118 7534 14170
rect 7714 14118 7716 14170
rect 7470 14116 7476 14118
rect 7532 14116 7556 14118
rect 7612 14116 7636 14118
rect 7692 14116 7716 14118
rect 7772 14116 7778 14118
rect 7470 14107 7778 14116
rect 12185 14172 12493 14181
rect 12185 14170 12191 14172
rect 12247 14170 12271 14172
rect 12327 14170 12351 14172
rect 12407 14170 12431 14172
rect 12487 14170 12493 14172
rect 12247 14118 12249 14170
rect 12429 14118 12431 14170
rect 12185 14116 12191 14118
rect 12247 14116 12271 14118
rect 12327 14116 12351 14118
rect 12407 14116 12431 14118
rect 12487 14116 12493 14118
rect 12185 14107 12493 14116
rect 16900 14172 17208 14181
rect 16900 14170 16906 14172
rect 16962 14170 16986 14172
rect 17042 14170 17066 14172
rect 17122 14170 17146 14172
rect 17202 14170 17208 14172
rect 16962 14118 16964 14170
rect 17144 14118 17146 14170
rect 16900 14116 16906 14118
rect 16962 14116 16986 14118
rect 17042 14116 17066 14118
rect 17122 14116 17146 14118
rect 17202 14116 17208 14118
rect 16900 14107 17208 14116
rect 5112 13628 5420 13637
rect 5112 13626 5118 13628
rect 5174 13626 5198 13628
rect 5254 13626 5278 13628
rect 5334 13626 5358 13628
rect 5414 13626 5420 13628
rect 5174 13574 5176 13626
rect 5356 13574 5358 13626
rect 5112 13572 5118 13574
rect 5174 13572 5198 13574
rect 5254 13572 5278 13574
rect 5334 13572 5358 13574
rect 5414 13572 5420 13574
rect 5112 13563 5420 13572
rect 9827 13628 10135 13637
rect 9827 13626 9833 13628
rect 9889 13626 9913 13628
rect 9969 13626 9993 13628
rect 10049 13626 10073 13628
rect 10129 13626 10135 13628
rect 9889 13574 9891 13626
rect 10071 13574 10073 13626
rect 9827 13572 9833 13574
rect 9889 13572 9913 13574
rect 9969 13572 9993 13574
rect 10049 13572 10073 13574
rect 10129 13572 10135 13574
rect 9827 13563 10135 13572
rect 14542 13628 14850 13637
rect 14542 13626 14548 13628
rect 14604 13626 14628 13628
rect 14684 13626 14708 13628
rect 14764 13626 14788 13628
rect 14844 13626 14850 13628
rect 14604 13574 14606 13626
rect 14786 13574 14788 13626
rect 14542 13572 14548 13574
rect 14604 13572 14628 13574
rect 14684 13572 14708 13574
rect 14764 13572 14788 13574
rect 14844 13572 14850 13574
rect 14542 13563 14850 13572
rect 19257 13628 19565 13637
rect 19257 13626 19263 13628
rect 19319 13626 19343 13628
rect 19399 13626 19423 13628
rect 19479 13626 19503 13628
rect 19559 13626 19565 13628
rect 19319 13574 19321 13626
rect 19501 13574 19503 13626
rect 19257 13572 19263 13574
rect 19319 13572 19343 13574
rect 19399 13572 19423 13574
rect 19479 13572 19503 13574
rect 19559 13572 19565 13574
rect 19257 13563 19565 13572
rect 2755 13084 3063 13093
rect 2755 13082 2761 13084
rect 2817 13082 2841 13084
rect 2897 13082 2921 13084
rect 2977 13082 3001 13084
rect 3057 13082 3063 13084
rect 2817 13030 2819 13082
rect 2999 13030 3001 13082
rect 2755 13028 2761 13030
rect 2817 13028 2841 13030
rect 2897 13028 2921 13030
rect 2977 13028 3001 13030
rect 3057 13028 3063 13030
rect 2755 13019 3063 13028
rect 7470 13084 7778 13093
rect 7470 13082 7476 13084
rect 7532 13082 7556 13084
rect 7612 13082 7636 13084
rect 7692 13082 7716 13084
rect 7772 13082 7778 13084
rect 7532 13030 7534 13082
rect 7714 13030 7716 13082
rect 7470 13028 7476 13030
rect 7532 13028 7556 13030
rect 7612 13028 7636 13030
rect 7692 13028 7716 13030
rect 7772 13028 7778 13030
rect 7470 13019 7778 13028
rect 12185 13084 12493 13093
rect 12185 13082 12191 13084
rect 12247 13082 12271 13084
rect 12327 13082 12351 13084
rect 12407 13082 12431 13084
rect 12487 13082 12493 13084
rect 12247 13030 12249 13082
rect 12429 13030 12431 13082
rect 12185 13028 12191 13030
rect 12247 13028 12271 13030
rect 12327 13028 12351 13030
rect 12407 13028 12431 13030
rect 12487 13028 12493 13030
rect 12185 13019 12493 13028
rect 16900 13084 17208 13093
rect 16900 13082 16906 13084
rect 16962 13082 16986 13084
rect 17042 13082 17066 13084
rect 17122 13082 17146 13084
rect 17202 13082 17208 13084
rect 16962 13030 16964 13082
rect 17144 13030 17146 13082
rect 16900 13028 16906 13030
rect 16962 13028 16986 13030
rect 17042 13028 17066 13030
rect 17122 13028 17146 13030
rect 17202 13028 17208 13030
rect 16900 13019 17208 13028
rect 5112 12540 5420 12549
rect 5112 12538 5118 12540
rect 5174 12538 5198 12540
rect 5254 12538 5278 12540
rect 5334 12538 5358 12540
rect 5414 12538 5420 12540
rect 5174 12486 5176 12538
rect 5356 12486 5358 12538
rect 5112 12484 5118 12486
rect 5174 12484 5198 12486
rect 5254 12484 5278 12486
rect 5334 12484 5358 12486
rect 5414 12484 5420 12486
rect 5112 12475 5420 12484
rect 9827 12540 10135 12549
rect 9827 12538 9833 12540
rect 9889 12538 9913 12540
rect 9969 12538 9993 12540
rect 10049 12538 10073 12540
rect 10129 12538 10135 12540
rect 9889 12486 9891 12538
rect 10071 12486 10073 12538
rect 9827 12484 9833 12486
rect 9889 12484 9913 12486
rect 9969 12484 9993 12486
rect 10049 12484 10073 12486
rect 10129 12484 10135 12486
rect 9827 12475 10135 12484
rect 14542 12540 14850 12549
rect 14542 12538 14548 12540
rect 14604 12538 14628 12540
rect 14684 12538 14708 12540
rect 14764 12538 14788 12540
rect 14844 12538 14850 12540
rect 14604 12486 14606 12538
rect 14786 12486 14788 12538
rect 14542 12484 14548 12486
rect 14604 12484 14628 12486
rect 14684 12484 14708 12486
rect 14764 12484 14788 12486
rect 14844 12484 14850 12486
rect 14542 12475 14850 12484
rect 19257 12540 19565 12549
rect 19257 12538 19263 12540
rect 19319 12538 19343 12540
rect 19399 12538 19423 12540
rect 19479 12538 19503 12540
rect 19559 12538 19565 12540
rect 19319 12486 19321 12538
rect 19501 12486 19503 12538
rect 19257 12484 19263 12486
rect 19319 12484 19343 12486
rect 19399 12484 19423 12486
rect 19479 12484 19503 12486
rect 19559 12484 19565 12486
rect 19257 12475 19565 12484
rect 2755 11996 3063 12005
rect 2755 11994 2761 11996
rect 2817 11994 2841 11996
rect 2897 11994 2921 11996
rect 2977 11994 3001 11996
rect 3057 11994 3063 11996
rect 2817 11942 2819 11994
rect 2999 11942 3001 11994
rect 2755 11940 2761 11942
rect 2817 11940 2841 11942
rect 2897 11940 2921 11942
rect 2977 11940 3001 11942
rect 3057 11940 3063 11942
rect 2755 11931 3063 11940
rect 7470 11996 7778 12005
rect 7470 11994 7476 11996
rect 7532 11994 7556 11996
rect 7612 11994 7636 11996
rect 7692 11994 7716 11996
rect 7772 11994 7778 11996
rect 7532 11942 7534 11994
rect 7714 11942 7716 11994
rect 7470 11940 7476 11942
rect 7532 11940 7556 11942
rect 7612 11940 7636 11942
rect 7692 11940 7716 11942
rect 7772 11940 7778 11942
rect 7470 11931 7778 11940
rect 12185 11996 12493 12005
rect 12185 11994 12191 11996
rect 12247 11994 12271 11996
rect 12327 11994 12351 11996
rect 12407 11994 12431 11996
rect 12487 11994 12493 11996
rect 12247 11942 12249 11994
rect 12429 11942 12431 11994
rect 12185 11940 12191 11942
rect 12247 11940 12271 11942
rect 12327 11940 12351 11942
rect 12407 11940 12431 11942
rect 12487 11940 12493 11942
rect 12185 11931 12493 11940
rect 16900 11996 17208 12005
rect 16900 11994 16906 11996
rect 16962 11994 16986 11996
rect 17042 11994 17066 11996
rect 17122 11994 17146 11996
rect 17202 11994 17208 11996
rect 16962 11942 16964 11994
rect 17144 11942 17146 11994
rect 16900 11940 16906 11942
rect 16962 11940 16986 11942
rect 17042 11940 17066 11942
rect 17122 11940 17146 11942
rect 17202 11940 17208 11942
rect 16900 11931 17208 11940
rect 5112 11452 5420 11461
rect 5112 11450 5118 11452
rect 5174 11450 5198 11452
rect 5254 11450 5278 11452
rect 5334 11450 5358 11452
rect 5414 11450 5420 11452
rect 5174 11398 5176 11450
rect 5356 11398 5358 11450
rect 5112 11396 5118 11398
rect 5174 11396 5198 11398
rect 5254 11396 5278 11398
rect 5334 11396 5358 11398
rect 5414 11396 5420 11398
rect 5112 11387 5420 11396
rect 9827 11452 10135 11461
rect 9827 11450 9833 11452
rect 9889 11450 9913 11452
rect 9969 11450 9993 11452
rect 10049 11450 10073 11452
rect 10129 11450 10135 11452
rect 9889 11398 9891 11450
rect 10071 11398 10073 11450
rect 9827 11396 9833 11398
rect 9889 11396 9913 11398
rect 9969 11396 9993 11398
rect 10049 11396 10073 11398
rect 10129 11396 10135 11398
rect 9827 11387 10135 11396
rect 14542 11452 14850 11461
rect 14542 11450 14548 11452
rect 14604 11450 14628 11452
rect 14684 11450 14708 11452
rect 14764 11450 14788 11452
rect 14844 11450 14850 11452
rect 14604 11398 14606 11450
rect 14786 11398 14788 11450
rect 14542 11396 14548 11398
rect 14604 11396 14628 11398
rect 14684 11396 14708 11398
rect 14764 11396 14788 11398
rect 14844 11396 14850 11398
rect 14542 11387 14850 11396
rect 19257 11452 19565 11461
rect 19257 11450 19263 11452
rect 19319 11450 19343 11452
rect 19399 11450 19423 11452
rect 19479 11450 19503 11452
rect 19559 11450 19565 11452
rect 19319 11398 19321 11450
rect 19501 11398 19503 11450
rect 19257 11396 19263 11398
rect 19319 11396 19343 11398
rect 19399 11396 19423 11398
rect 19479 11396 19503 11398
rect 19559 11396 19565 11398
rect 19257 11387 19565 11396
rect 2755 10908 3063 10917
rect 2755 10906 2761 10908
rect 2817 10906 2841 10908
rect 2897 10906 2921 10908
rect 2977 10906 3001 10908
rect 3057 10906 3063 10908
rect 2817 10854 2819 10906
rect 2999 10854 3001 10906
rect 2755 10852 2761 10854
rect 2817 10852 2841 10854
rect 2897 10852 2921 10854
rect 2977 10852 3001 10854
rect 3057 10852 3063 10854
rect 2755 10843 3063 10852
rect 7470 10908 7778 10917
rect 7470 10906 7476 10908
rect 7532 10906 7556 10908
rect 7612 10906 7636 10908
rect 7692 10906 7716 10908
rect 7772 10906 7778 10908
rect 7532 10854 7534 10906
rect 7714 10854 7716 10906
rect 7470 10852 7476 10854
rect 7532 10852 7556 10854
rect 7612 10852 7636 10854
rect 7692 10852 7716 10854
rect 7772 10852 7778 10854
rect 7470 10843 7778 10852
rect 12185 10908 12493 10917
rect 12185 10906 12191 10908
rect 12247 10906 12271 10908
rect 12327 10906 12351 10908
rect 12407 10906 12431 10908
rect 12487 10906 12493 10908
rect 12247 10854 12249 10906
rect 12429 10854 12431 10906
rect 12185 10852 12191 10854
rect 12247 10852 12271 10854
rect 12327 10852 12351 10854
rect 12407 10852 12431 10854
rect 12487 10852 12493 10854
rect 12185 10843 12493 10852
rect 16900 10908 17208 10917
rect 16900 10906 16906 10908
rect 16962 10906 16986 10908
rect 17042 10906 17066 10908
rect 17122 10906 17146 10908
rect 17202 10906 17208 10908
rect 16962 10854 16964 10906
rect 17144 10854 17146 10906
rect 16900 10852 16906 10854
rect 16962 10852 16986 10854
rect 17042 10852 17066 10854
rect 17122 10852 17146 10854
rect 17202 10852 17208 10854
rect 16900 10843 17208 10852
rect 5112 10364 5420 10373
rect 5112 10362 5118 10364
rect 5174 10362 5198 10364
rect 5254 10362 5278 10364
rect 5334 10362 5358 10364
rect 5414 10362 5420 10364
rect 5174 10310 5176 10362
rect 5356 10310 5358 10362
rect 5112 10308 5118 10310
rect 5174 10308 5198 10310
rect 5254 10308 5278 10310
rect 5334 10308 5358 10310
rect 5414 10308 5420 10310
rect 5112 10299 5420 10308
rect 9827 10364 10135 10373
rect 9827 10362 9833 10364
rect 9889 10362 9913 10364
rect 9969 10362 9993 10364
rect 10049 10362 10073 10364
rect 10129 10362 10135 10364
rect 9889 10310 9891 10362
rect 10071 10310 10073 10362
rect 9827 10308 9833 10310
rect 9889 10308 9913 10310
rect 9969 10308 9993 10310
rect 10049 10308 10073 10310
rect 10129 10308 10135 10310
rect 9827 10299 10135 10308
rect 14542 10364 14850 10373
rect 14542 10362 14548 10364
rect 14604 10362 14628 10364
rect 14684 10362 14708 10364
rect 14764 10362 14788 10364
rect 14844 10362 14850 10364
rect 14604 10310 14606 10362
rect 14786 10310 14788 10362
rect 14542 10308 14548 10310
rect 14604 10308 14628 10310
rect 14684 10308 14708 10310
rect 14764 10308 14788 10310
rect 14844 10308 14850 10310
rect 14542 10299 14850 10308
rect 19257 10364 19565 10373
rect 19257 10362 19263 10364
rect 19319 10362 19343 10364
rect 19399 10362 19423 10364
rect 19479 10362 19503 10364
rect 19559 10362 19565 10364
rect 19319 10310 19321 10362
rect 19501 10310 19503 10362
rect 19257 10308 19263 10310
rect 19319 10308 19343 10310
rect 19399 10308 19423 10310
rect 19479 10308 19503 10310
rect 19559 10308 19565 10310
rect 19257 10299 19565 10308
rect 19064 9920 19116 9926
rect 19062 9888 19064 9897
rect 19116 9888 19118 9897
rect 2755 9820 3063 9829
rect 2755 9818 2761 9820
rect 2817 9818 2841 9820
rect 2897 9818 2921 9820
rect 2977 9818 3001 9820
rect 3057 9818 3063 9820
rect 2817 9766 2819 9818
rect 2999 9766 3001 9818
rect 2755 9764 2761 9766
rect 2817 9764 2841 9766
rect 2897 9764 2921 9766
rect 2977 9764 3001 9766
rect 3057 9764 3063 9766
rect 2755 9755 3063 9764
rect 7470 9820 7778 9829
rect 7470 9818 7476 9820
rect 7532 9818 7556 9820
rect 7612 9818 7636 9820
rect 7692 9818 7716 9820
rect 7772 9818 7778 9820
rect 7532 9766 7534 9818
rect 7714 9766 7716 9818
rect 7470 9764 7476 9766
rect 7532 9764 7556 9766
rect 7612 9764 7636 9766
rect 7692 9764 7716 9766
rect 7772 9764 7778 9766
rect 7470 9755 7778 9764
rect 12185 9820 12493 9829
rect 12185 9818 12191 9820
rect 12247 9818 12271 9820
rect 12327 9818 12351 9820
rect 12407 9818 12431 9820
rect 12487 9818 12493 9820
rect 12247 9766 12249 9818
rect 12429 9766 12431 9818
rect 12185 9764 12191 9766
rect 12247 9764 12271 9766
rect 12327 9764 12351 9766
rect 12407 9764 12431 9766
rect 12487 9764 12493 9766
rect 12185 9755 12493 9764
rect 16900 9820 17208 9829
rect 19062 9823 19118 9832
rect 16900 9818 16906 9820
rect 16962 9818 16986 9820
rect 17042 9818 17066 9820
rect 17122 9818 17146 9820
rect 17202 9818 17208 9820
rect 16962 9766 16964 9818
rect 17144 9766 17146 9818
rect 16900 9764 16906 9766
rect 16962 9764 16986 9766
rect 17042 9764 17066 9766
rect 17122 9764 17146 9766
rect 17202 9764 17208 9766
rect 16900 9755 17208 9764
rect 5112 9276 5420 9285
rect 5112 9274 5118 9276
rect 5174 9274 5198 9276
rect 5254 9274 5278 9276
rect 5334 9274 5358 9276
rect 5414 9274 5420 9276
rect 5174 9222 5176 9274
rect 5356 9222 5358 9274
rect 5112 9220 5118 9222
rect 5174 9220 5198 9222
rect 5254 9220 5278 9222
rect 5334 9220 5358 9222
rect 5414 9220 5420 9222
rect 5112 9211 5420 9220
rect 9827 9276 10135 9285
rect 9827 9274 9833 9276
rect 9889 9274 9913 9276
rect 9969 9274 9993 9276
rect 10049 9274 10073 9276
rect 10129 9274 10135 9276
rect 9889 9222 9891 9274
rect 10071 9222 10073 9274
rect 9827 9220 9833 9222
rect 9889 9220 9913 9222
rect 9969 9220 9993 9222
rect 10049 9220 10073 9222
rect 10129 9220 10135 9222
rect 9827 9211 10135 9220
rect 14542 9276 14850 9285
rect 14542 9274 14548 9276
rect 14604 9274 14628 9276
rect 14684 9274 14708 9276
rect 14764 9274 14788 9276
rect 14844 9274 14850 9276
rect 14604 9222 14606 9274
rect 14786 9222 14788 9274
rect 14542 9220 14548 9222
rect 14604 9220 14628 9222
rect 14684 9220 14708 9222
rect 14764 9220 14788 9222
rect 14844 9220 14850 9222
rect 14542 9211 14850 9220
rect 19257 9276 19565 9285
rect 19257 9274 19263 9276
rect 19319 9274 19343 9276
rect 19399 9274 19423 9276
rect 19479 9274 19503 9276
rect 19559 9274 19565 9276
rect 19319 9222 19321 9274
rect 19501 9222 19503 9274
rect 19257 9220 19263 9222
rect 19319 9220 19343 9222
rect 19399 9220 19423 9222
rect 19479 9220 19503 9222
rect 19559 9220 19565 9222
rect 19257 9211 19565 9220
rect 2755 8732 3063 8741
rect 2755 8730 2761 8732
rect 2817 8730 2841 8732
rect 2897 8730 2921 8732
rect 2977 8730 3001 8732
rect 3057 8730 3063 8732
rect 2817 8678 2819 8730
rect 2999 8678 3001 8730
rect 2755 8676 2761 8678
rect 2817 8676 2841 8678
rect 2897 8676 2921 8678
rect 2977 8676 3001 8678
rect 3057 8676 3063 8678
rect 2755 8667 3063 8676
rect 7470 8732 7778 8741
rect 7470 8730 7476 8732
rect 7532 8730 7556 8732
rect 7612 8730 7636 8732
rect 7692 8730 7716 8732
rect 7772 8730 7778 8732
rect 7532 8678 7534 8730
rect 7714 8678 7716 8730
rect 7470 8676 7476 8678
rect 7532 8676 7556 8678
rect 7612 8676 7636 8678
rect 7692 8676 7716 8678
rect 7772 8676 7778 8678
rect 7470 8667 7778 8676
rect 12185 8732 12493 8741
rect 12185 8730 12191 8732
rect 12247 8730 12271 8732
rect 12327 8730 12351 8732
rect 12407 8730 12431 8732
rect 12487 8730 12493 8732
rect 12247 8678 12249 8730
rect 12429 8678 12431 8730
rect 12185 8676 12191 8678
rect 12247 8676 12271 8678
rect 12327 8676 12351 8678
rect 12407 8676 12431 8678
rect 12487 8676 12493 8678
rect 12185 8667 12493 8676
rect 16900 8732 17208 8741
rect 16900 8730 16906 8732
rect 16962 8730 16986 8732
rect 17042 8730 17066 8732
rect 17122 8730 17146 8732
rect 17202 8730 17208 8732
rect 16962 8678 16964 8730
rect 17144 8678 17146 8730
rect 16900 8676 16906 8678
rect 16962 8676 16986 8678
rect 17042 8676 17066 8678
rect 17122 8676 17146 8678
rect 17202 8676 17208 8678
rect 16900 8667 17208 8676
rect 5112 8188 5420 8197
rect 5112 8186 5118 8188
rect 5174 8186 5198 8188
rect 5254 8186 5278 8188
rect 5334 8186 5358 8188
rect 5414 8186 5420 8188
rect 5174 8134 5176 8186
rect 5356 8134 5358 8186
rect 5112 8132 5118 8134
rect 5174 8132 5198 8134
rect 5254 8132 5278 8134
rect 5334 8132 5358 8134
rect 5414 8132 5420 8134
rect 5112 8123 5420 8132
rect 9827 8188 10135 8197
rect 9827 8186 9833 8188
rect 9889 8186 9913 8188
rect 9969 8186 9993 8188
rect 10049 8186 10073 8188
rect 10129 8186 10135 8188
rect 9889 8134 9891 8186
rect 10071 8134 10073 8186
rect 9827 8132 9833 8134
rect 9889 8132 9913 8134
rect 9969 8132 9993 8134
rect 10049 8132 10073 8134
rect 10129 8132 10135 8134
rect 9827 8123 10135 8132
rect 14542 8188 14850 8197
rect 14542 8186 14548 8188
rect 14604 8186 14628 8188
rect 14684 8186 14708 8188
rect 14764 8186 14788 8188
rect 14844 8186 14850 8188
rect 14604 8134 14606 8186
rect 14786 8134 14788 8186
rect 14542 8132 14548 8134
rect 14604 8132 14628 8134
rect 14684 8132 14708 8134
rect 14764 8132 14788 8134
rect 14844 8132 14850 8134
rect 14542 8123 14850 8132
rect 19257 8188 19565 8197
rect 19257 8186 19263 8188
rect 19319 8186 19343 8188
rect 19399 8186 19423 8188
rect 19479 8186 19503 8188
rect 19559 8186 19565 8188
rect 19319 8134 19321 8186
rect 19501 8134 19503 8186
rect 19257 8132 19263 8134
rect 19319 8132 19343 8134
rect 19399 8132 19423 8134
rect 19479 8132 19503 8134
rect 19559 8132 19565 8134
rect 19257 8123 19565 8132
rect 2755 7644 3063 7653
rect 2755 7642 2761 7644
rect 2817 7642 2841 7644
rect 2897 7642 2921 7644
rect 2977 7642 3001 7644
rect 3057 7642 3063 7644
rect 2817 7590 2819 7642
rect 2999 7590 3001 7642
rect 2755 7588 2761 7590
rect 2817 7588 2841 7590
rect 2897 7588 2921 7590
rect 2977 7588 3001 7590
rect 3057 7588 3063 7590
rect 2755 7579 3063 7588
rect 7470 7644 7778 7653
rect 7470 7642 7476 7644
rect 7532 7642 7556 7644
rect 7612 7642 7636 7644
rect 7692 7642 7716 7644
rect 7772 7642 7778 7644
rect 7532 7590 7534 7642
rect 7714 7590 7716 7642
rect 7470 7588 7476 7590
rect 7532 7588 7556 7590
rect 7612 7588 7636 7590
rect 7692 7588 7716 7590
rect 7772 7588 7778 7590
rect 7470 7579 7778 7588
rect 12185 7644 12493 7653
rect 12185 7642 12191 7644
rect 12247 7642 12271 7644
rect 12327 7642 12351 7644
rect 12407 7642 12431 7644
rect 12487 7642 12493 7644
rect 12247 7590 12249 7642
rect 12429 7590 12431 7642
rect 12185 7588 12191 7590
rect 12247 7588 12271 7590
rect 12327 7588 12351 7590
rect 12407 7588 12431 7590
rect 12487 7588 12493 7590
rect 12185 7579 12493 7588
rect 16900 7644 17208 7653
rect 16900 7642 16906 7644
rect 16962 7642 16986 7644
rect 17042 7642 17066 7644
rect 17122 7642 17146 7644
rect 17202 7642 17208 7644
rect 16962 7590 16964 7642
rect 17144 7590 17146 7642
rect 16900 7588 16906 7590
rect 16962 7588 16986 7590
rect 17042 7588 17066 7590
rect 17122 7588 17146 7590
rect 17202 7588 17208 7590
rect 16900 7579 17208 7588
rect 5112 7100 5420 7109
rect 5112 7098 5118 7100
rect 5174 7098 5198 7100
rect 5254 7098 5278 7100
rect 5334 7098 5358 7100
rect 5414 7098 5420 7100
rect 5174 7046 5176 7098
rect 5356 7046 5358 7098
rect 5112 7044 5118 7046
rect 5174 7044 5198 7046
rect 5254 7044 5278 7046
rect 5334 7044 5358 7046
rect 5414 7044 5420 7046
rect 5112 7035 5420 7044
rect 9827 7100 10135 7109
rect 9827 7098 9833 7100
rect 9889 7098 9913 7100
rect 9969 7098 9993 7100
rect 10049 7098 10073 7100
rect 10129 7098 10135 7100
rect 9889 7046 9891 7098
rect 10071 7046 10073 7098
rect 9827 7044 9833 7046
rect 9889 7044 9913 7046
rect 9969 7044 9993 7046
rect 10049 7044 10073 7046
rect 10129 7044 10135 7046
rect 9827 7035 10135 7044
rect 14542 7100 14850 7109
rect 14542 7098 14548 7100
rect 14604 7098 14628 7100
rect 14684 7098 14708 7100
rect 14764 7098 14788 7100
rect 14844 7098 14850 7100
rect 14604 7046 14606 7098
rect 14786 7046 14788 7098
rect 14542 7044 14548 7046
rect 14604 7044 14628 7046
rect 14684 7044 14708 7046
rect 14764 7044 14788 7046
rect 14844 7044 14850 7046
rect 14542 7035 14850 7044
rect 19257 7100 19565 7109
rect 19257 7098 19263 7100
rect 19319 7098 19343 7100
rect 19399 7098 19423 7100
rect 19479 7098 19503 7100
rect 19559 7098 19565 7100
rect 19319 7046 19321 7098
rect 19501 7046 19503 7098
rect 19257 7044 19263 7046
rect 19319 7044 19343 7046
rect 19399 7044 19423 7046
rect 19479 7044 19503 7046
rect 19559 7044 19565 7046
rect 19257 7035 19565 7044
rect 2755 6556 3063 6565
rect 2755 6554 2761 6556
rect 2817 6554 2841 6556
rect 2897 6554 2921 6556
rect 2977 6554 3001 6556
rect 3057 6554 3063 6556
rect 2817 6502 2819 6554
rect 2999 6502 3001 6554
rect 2755 6500 2761 6502
rect 2817 6500 2841 6502
rect 2897 6500 2921 6502
rect 2977 6500 3001 6502
rect 3057 6500 3063 6502
rect 2755 6491 3063 6500
rect 7470 6556 7778 6565
rect 7470 6554 7476 6556
rect 7532 6554 7556 6556
rect 7612 6554 7636 6556
rect 7692 6554 7716 6556
rect 7772 6554 7778 6556
rect 7532 6502 7534 6554
rect 7714 6502 7716 6554
rect 7470 6500 7476 6502
rect 7532 6500 7556 6502
rect 7612 6500 7636 6502
rect 7692 6500 7716 6502
rect 7772 6500 7778 6502
rect 7470 6491 7778 6500
rect 12185 6556 12493 6565
rect 12185 6554 12191 6556
rect 12247 6554 12271 6556
rect 12327 6554 12351 6556
rect 12407 6554 12431 6556
rect 12487 6554 12493 6556
rect 12247 6502 12249 6554
rect 12429 6502 12431 6554
rect 12185 6500 12191 6502
rect 12247 6500 12271 6502
rect 12327 6500 12351 6502
rect 12407 6500 12431 6502
rect 12487 6500 12493 6502
rect 12185 6491 12493 6500
rect 16900 6556 17208 6565
rect 16900 6554 16906 6556
rect 16962 6554 16986 6556
rect 17042 6554 17066 6556
rect 17122 6554 17146 6556
rect 17202 6554 17208 6556
rect 16962 6502 16964 6554
rect 17144 6502 17146 6554
rect 16900 6500 16906 6502
rect 16962 6500 16986 6502
rect 17042 6500 17066 6502
rect 17122 6500 17146 6502
rect 17202 6500 17208 6502
rect 16900 6491 17208 6500
rect 5112 6012 5420 6021
rect 5112 6010 5118 6012
rect 5174 6010 5198 6012
rect 5254 6010 5278 6012
rect 5334 6010 5358 6012
rect 5414 6010 5420 6012
rect 5174 5958 5176 6010
rect 5356 5958 5358 6010
rect 5112 5956 5118 5958
rect 5174 5956 5198 5958
rect 5254 5956 5278 5958
rect 5334 5956 5358 5958
rect 5414 5956 5420 5958
rect 5112 5947 5420 5956
rect 9827 6012 10135 6021
rect 9827 6010 9833 6012
rect 9889 6010 9913 6012
rect 9969 6010 9993 6012
rect 10049 6010 10073 6012
rect 10129 6010 10135 6012
rect 9889 5958 9891 6010
rect 10071 5958 10073 6010
rect 9827 5956 9833 5958
rect 9889 5956 9913 5958
rect 9969 5956 9993 5958
rect 10049 5956 10073 5958
rect 10129 5956 10135 5958
rect 9827 5947 10135 5956
rect 14542 6012 14850 6021
rect 14542 6010 14548 6012
rect 14604 6010 14628 6012
rect 14684 6010 14708 6012
rect 14764 6010 14788 6012
rect 14844 6010 14850 6012
rect 14604 5958 14606 6010
rect 14786 5958 14788 6010
rect 14542 5956 14548 5958
rect 14604 5956 14628 5958
rect 14684 5956 14708 5958
rect 14764 5956 14788 5958
rect 14844 5956 14850 5958
rect 14542 5947 14850 5956
rect 19257 6012 19565 6021
rect 19257 6010 19263 6012
rect 19319 6010 19343 6012
rect 19399 6010 19423 6012
rect 19479 6010 19503 6012
rect 19559 6010 19565 6012
rect 19319 5958 19321 6010
rect 19501 5958 19503 6010
rect 19257 5956 19263 5958
rect 19319 5956 19343 5958
rect 19399 5956 19423 5958
rect 19479 5956 19503 5958
rect 19559 5956 19565 5958
rect 19257 5947 19565 5956
rect 2755 5468 3063 5477
rect 2755 5466 2761 5468
rect 2817 5466 2841 5468
rect 2897 5466 2921 5468
rect 2977 5466 3001 5468
rect 3057 5466 3063 5468
rect 2817 5414 2819 5466
rect 2999 5414 3001 5466
rect 2755 5412 2761 5414
rect 2817 5412 2841 5414
rect 2897 5412 2921 5414
rect 2977 5412 3001 5414
rect 3057 5412 3063 5414
rect 2755 5403 3063 5412
rect 7470 5468 7778 5477
rect 7470 5466 7476 5468
rect 7532 5466 7556 5468
rect 7612 5466 7636 5468
rect 7692 5466 7716 5468
rect 7772 5466 7778 5468
rect 7532 5414 7534 5466
rect 7714 5414 7716 5466
rect 7470 5412 7476 5414
rect 7532 5412 7556 5414
rect 7612 5412 7636 5414
rect 7692 5412 7716 5414
rect 7772 5412 7778 5414
rect 7470 5403 7778 5412
rect 12185 5468 12493 5477
rect 12185 5466 12191 5468
rect 12247 5466 12271 5468
rect 12327 5466 12351 5468
rect 12407 5466 12431 5468
rect 12487 5466 12493 5468
rect 12247 5414 12249 5466
rect 12429 5414 12431 5466
rect 12185 5412 12191 5414
rect 12247 5412 12271 5414
rect 12327 5412 12351 5414
rect 12407 5412 12431 5414
rect 12487 5412 12493 5414
rect 12185 5403 12493 5412
rect 16900 5468 17208 5477
rect 16900 5466 16906 5468
rect 16962 5466 16986 5468
rect 17042 5466 17066 5468
rect 17122 5466 17146 5468
rect 17202 5466 17208 5468
rect 16962 5414 16964 5466
rect 17144 5414 17146 5466
rect 16900 5412 16906 5414
rect 16962 5412 16986 5414
rect 17042 5412 17066 5414
rect 17122 5412 17146 5414
rect 17202 5412 17208 5414
rect 16900 5403 17208 5412
rect 5112 4924 5420 4933
rect 5112 4922 5118 4924
rect 5174 4922 5198 4924
rect 5254 4922 5278 4924
rect 5334 4922 5358 4924
rect 5414 4922 5420 4924
rect 5174 4870 5176 4922
rect 5356 4870 5358 4922
rect 5112 4868 5118 4870
rect 5174 4868 5198 4870
rect 5254 4868 5278 4870
rect 5334 4868 5358 4870
rect 5414 4868 5420 4870
rect 5112 4859 5420 4868
rect 9827 4924 10135 4933
rect 9827 4922 9833 4924
rect 9889 4922 9913 4924
rect 9969 4922 9993 4924
rect 10049 4922 10073 4924
rect 10129 4922 10135 4924
rect 9889 4870 9891 4922
rect 10071 4870 10073 4922
rect 9827 4868 9833 4870
rect 9889 4868 9913 4870
rect 9969 4868 9993 4870
rect 10049 4868 10073 4870
rect 10129 4868 10135 4870
rect 9827 4859 10135 4868
rect 14542 4924 14850 4933
rect 14542 4922 14548 4924
rect 14604 4922 14628 4924
rect 14684 4922 14708 4924
rect 14764 4922 14788 4924
rect 14844 4922 14850 4924
rect 14604 4870 14606 4922
rect 14786 4870 14788 4922
rect 14542 4868 14548 4870
rect 14604 4868 14628 4870
rect 14684 4868 14708 4870
rect 14764 4868 14788 4870
rect 14844 4868 14850 4870
rect 14542 4859 14850 4868
rect 19257 4924 19565 4933
rect 19257 4922 19263 4924
rect 19319 4922 19343 4924
rect 19399 4922 19423 4924
rect 19479 4922 19503 4924
rect 19559 4922 19565 4924
rect 19319 4870 19321 4922
rect 19501 4870 19503 4922
rect 19257 4868 19263 4870
rect 19319 4868 19343 4870
rect 19399 4868 19423 4870
rect 19479 4868 19503 4870
rect 19559 4868 19565 4870
rect 19257 4859 19565 4868
rect 2755 4380 3063 4389
rect 2755 4378 2761 4380
rect 2817 4378 2841 4380
rect 2897 4378 2921 4380
rect 2977 4378 3001 4380
rect 3057 4378 3063 4380
rect 2817 4326 2819 4378
rect 2999 4326 3001 4378
rect 2755 4324 2761 4326
rect 2817 4324 2841 4326
rect 2897 4324 2921 4326
rect 2977 4324 3001 4326
rect 3057 4324 3063 4326
rect 2755 4315 3063 4324
rect 7470 4380 7778 4389
rect 7470 4378 7476 4380
rect 7532 4378 7556 4380
rect 7612 4378 7636 4380
rect 7692 4378 7716 4380
rect 7772 4378 7778 4380
rect 7532 4326 7534 4378
rect 7714 4326 7716 4378
rect 7470 4324 7476 4326
rect 7532 4324 7556 4326
rect 7612 4324 7636 4326
rect 7692 4324 7716 4326
rect 7772 4324 7778 4326
rect 7470 4315 7778 4324
rect 12185 4380 12493 4389
rect 12185 4378 12191 4380
rect 12247 4378 12271 4380
rect 12327 4378 12351 4380
rect 12407 4378 12431 4380
rect 12487 4378 12493 4380
rect 12247 4326 12249 4378
rect 12429 4326 12431 4378
rect 12185 4324 12191 4326
rect 12247 4324 12271 4326
rect 12327 4324 12351 4326
rect 12407 4324 12431 4326
rect 12487 4324 12493 4326
rect 12185 4315 12493 4324
rect 16900 4380 17208 4389
rect 16900 4378 16906 4380
rect 16962 4378 16986 4380
rect 17042 4378 17066 4380
rect 17122 4378 17146 4380
rect 17202 4378 17208 4380
rect 16962 4326 16964 4378
rect 17144 4326 17146 4378
rect 16900 4324 16906 4326
rect 16962 4324 16986 4326
rect 17042 4324 17066 4326
rect 17122 4324 17146 4326
rect 17202 4324 17208 4326
rect 16900 4315 17208 4324
rect 5112 3836 5420 3845
rect 5112 3834 5118 3836
rect 5174 3834 5198 3836
rect 5254 3834 5278 3836
rect 5334 3834 5358 3836
rect 5414 3834 5420 3836
rect 5174 3782 5176 3834
rect 5356 3782 5358 3834
rect 5112 3780 5118 3782
rect 5174 3780 5198 3782
rect 5254 3780 5278 3782
rect 5334 3780 5358 3782
rect 5414 3780 5420 3782
rect 5112 3771 5420 3780
rect 9827 3836 10135 3845
rect 9827 3834 9833 3836
rect 9889 3834 9913 3836
rect 9969 3834 9993 3836
rect 10049 3834 10073 3836
rect 10129 3834 10135 3836
rect 9889 3782 9891 3834
rect 10071 3782 10073 3834
rect 9827 3780 9833 3782
rect 9889 3780 9913 3782
rect 9969 3780 9993 3782
rect 10049 3780 10073 3782
rect 10129 3780 10135 3782
rect 9827 3771 10135 3780
rect 14542 3836 14850 3845
rect 14542 3834 14548 3836
rect 14604 3834 14628 3836
rect 14684 3834 14708 3836
rect 14764 3834 14788 3836
rect 14844 3834 14850 3836
rect 14604 3782 14606 3834
rect 14786 3782 14788 3834
rect 14542 3780 14548 3782
rect 14604 3780 14628 3782
rect 14684 3780 14708 3782
rect 14764 3780 14788 3782
rect 14844 3780 14850 3782
rect 14542 3771 14850 3780
rect 19257 3836 19565 3845
rect 19257 3834 19263 3836
rect 19319 3834 19343 3836
rect 19399 3834 19423 3836
rect 19479 3834 19503 3836
rect 19559 3834 19565 3836
rect 19319 3782 19321 3834
rect 19501 3782 19503 3834
rect 19257 3780 19263 3782
rect 19319 3780 19343 3782
rect 19399 3780 19423 3782
rect 19479 3780 19503 3782
rect 19559 3780 19565 3782
rect 19257 3771 19565 3780
rect 2755 3292 3063 3301
rect 2755 3290 2761 3292
rect 2817 3290 2841 3292
rect 2897 3290 2921 3292
rect 2977 3290 3001 3292
rect 3057 3290 3063 3292
rect 2817 3238 2819 3290
rect 2999 3238 3001 3290
rect 2755 3236 2761 3238
rect 2817 3236 2841 3238
rect 2897 3236 2921 3238
rect 2977 3236 3001 3238
rect 3057 3236 3063 3238
rect 2755 3227 3063 3236
rect 7470 3292 7778 3301
rect 7470 3290 7476 3292
rect 7532 3290 7556 3292
rect 7612 3290 7636 3292
rect 7692 3290 7716 3292
rect 7772 3290 7778 3292
rect 7532 3238 7534 3290
rect 7714 3238 7716 3290
rect 7470 3236 7476 3238
rect 7532 3236 7556 3238
rect 7612 3236 7636 3238
rect 7692 3236 7716 3238
rect 7772 3236 7778 3238
rect 7470 3227 7778 3236
rect 12185 3292 12493 3301
rect 12185 3290 12191 3292
rect 12247 3290 12271 3292
rect 12327 3290 12351 3292
rect 12407 3290 12431 3292
rect 12487 3290 12493 3292
rect 12247 3238 12249 3290
rect 12429 3238 12431 3290
rect 12185 3236 12191 3238
rect 12247 3236 12271 3238
rect 12327 3236 12351 3238
rect 12407 3236 12431 3238
rect 12487 3236 12493 3238
rect 12185 3227 12493 3236
rect 16900 3292 17208 3301
rect 16900 3290 16906 3292
rect 16962 3290 16986 3292
rect 17042 3290 17066 3292
rect 17122 3290 17146 3292
rect 17202 3290 17208 3292
rect 16962 3238 16964 3290
rect 17144 3238 17146 3290
rect 16900 3236 16906 3238
rect 16962 3236 16986 3238
rect 17042 3236 17066 3238
rect 17122 3236 17146 3238
rect 17202 3236 17208 3238
rect 16900 3227 17208 3236
rect 5112 2748 5420 2757
rect 5112 2746 5118 2748
rect 5174 2746 5198 2748
rect 5254 2746 5278 2748
rect 5334 2746 5358 2748
rect 5414 2746 5420 2748
rect 5174 2694 5176 2746
rect 5356 2694 5358 2746
rect 5112 2692 5118 2694
rect 5174 2692 5198 2694
rect 5254 2692 5278 2694
rect 5334 2692 5358 2694
rect 5414 2692 5420 2694
rect 5112 2683 5420 2692
rect 9827 2748 10135 2757
rect 9827 2746 9833 2748
rect 9889 2746 9913 2748
rect 9969 2746 9993 2748
rect 10049 2746 10073 2748
rect 10129 2746 10135 2748
rect 9889 2694 9891 2746
rect 10071 2694 10073 2746
rect 9827 2692 9833 2694
rect 9889 2692 9913 2694
rect 9969 2692 9993 2694
rect 10049 2692 10073 2694
rect 10129 2692 10135 2694
rect 9827 2683 10135 2692
rect 14542 2748 14850 2757
rect 14542 2746 14548 2748
rect 14604 2746 14628 2748
rect 14684 2746 14708 2748
rect 14764 2746 14788 2748
rect 14844 2746 14850 2748
rect 14604 2694 14606 2746
rect 14786 2694 14788 2746
rect 14542 2692 14548 2694
rect 14604 2692 14628 2694
rect 14684 2692 14708 2694
rect 14764 2692 14788 2694
rect 14844 2692 14850 2694
rect 14542 2683 14850 2692
rect 19257 2748 19565 2757
rect 19257 2746 19263 2748
rect 19319 2746 19343 2748
rect 19399 2746 19423 2748
rect 19479 2746 19503 2748
rect 19559 2746 19565 2748
rect 19319 2694 19321 2746
rect 19501 2694 19503 2746
rect 19257 2692 19263 2694
rect 19319 2692 19343 2694
rect 19399 2692 19423 2694
rect 19479 2692 19503 2694
rect 19559 2692 19565 2694
rect 19257 2683 19565 2692
rect 2755 2204 3063 2213
rect 2755 2202 2761 2204
rect 2817 2202 2841 2204
rect 2897 2202 2921 2204
rect 2977 2202 3001 2204
rect 3057 2202 3063 2204
rect 2817 2150 2819 2202
rect 2999 2150 3001 2202
rect 2755 2148 2761 2150
rect 2817 2148 2841 2150
rect 2897 2148 2921 2150
rect 2977 2148 3001 2150
rect 3057 2148 3063 2150
rect 2755 2139 3063 2148
rect 7470 2204 7778 2213
rect 7470 2202 7476 2204
rect 7532 2202 7556 2204
rect 7612 2202 7636 2204
rect 7692 2202 7716 2204
rect 7772 2202 7778 2204
rect 7532 2150 7534 2202
rect 7714 2150 7716 2202
rect 7470 2148 7476 2150
rect 7532 2148 7556 2150
rect 7612 2148 7636 2150
rect 7692 2148 7716 2150
rect 7772 2148 7778 2150
rect 7470 2139 7778 2148
rect 12185 2204 12493 2213
rect 12185 2202 12191 2204
rect 12247 2202 12271 2204
rect 12327 2202 12351 2204
rect 12407 2202 12431 2204
rect 12487 2202 12493 2204
rect 12247 2150 12249 2202
rect 12429 2150 12431 2202
rect 12185 2148 12191 2150
rect 12247 2148 12271 2150
rect 12327 2148 12351 2150
rect 12407 2148 12431 2150
rect 12487 2148 12493 2150
rect 12185 2139 12493 2148
rect 16900 2204 17208 2213
rect 16900 2202 16906 2204
rect 16962 2202 16986 2204
rect 17042 2202 17066 2204
rect 17122 2202 17146 2204
rect 17202 2202 17208 2204
rect 16962 2150 16964 2202
rect 17144 2150 17146 2202
rect 16900 2148 16906 2150
rect 16962 2148 16986 2150
rect 17042 2148 17066 2150
rect 17122 2148 17146 2150
rect 17202 2148 17208 2150
rect 16900 2139 17208 2148
rect 5112 1660 5420 1669
rect 5112 1658 5118 1660
rect 5174 1658 5198 1660
rect 5254 1658 5278 1660
rect 5334 1658 5358 1660
rect 5414 1658 5420 1660
rect 5174 1606 5176 1658
rect 5356 1606 5358 1658
rect 5112 1604 5118 1606
rect 5174 1604 5198 1606
rect 5254 1604 5278 1606
rect 5334 1604 5358 1606
rect 5414 1604 5420 1606
rect 5112 1595 5420 1604
rect 9827 1660 10135 1669
rect 9827 1658 9833 1660
rect 9889 1658 9913 1660
rect 9969 1658 9993 1660
rect 10049 1658 10073 1660
rect 10129 1658 10135 1660
rect 9889 1606 9891 1658
rect 10071 1606 10073 1658
rect 9827 1604 9833 1606
rect 9889 1604 9913 1606
rect 9969 1604 9993 1606
rect 10049 1604 10073 1606
rect 10129 1604 10135 1606
rect 9827 1595 10135 1604
rect 14542 1660 14850 1669
rect 14542 1658 14548 1660
rect 14604 1658 14628 1660
rect 14684 1658 14708 1660
rect 14764 1658 14788 1660
rect 14844 1658 14850 1660
rect 14604 1606 14606 1658
rect 14786 1606 14788 1658
rect 14542 1604 14548 1606
rect 14604 1604 14628 1606
rect 14684 1604 14708 1606
rect 14764 1604 14788 1606
rect 14844 1604 14850 1606
rect 14542 1595 14850 1604
rect 19257 1660 19565 1669
rect 19257 1658 19263 1660
rect 19319 1658 19343 1660
rect 19399 1658 19423 1660
rect 19479 1658 19503 1660
rect 19559 1658 19565 1660
rect 19319 1606 19321 1658
rect 19501 1606 19503 1658
rect 19257 1604 19263 1606
rect 19319 1604 19343 1606
rect 19399 1604 19423 1606
rect 19479 1604 19503 1606
rect 19559 1604 19565 1606
rect 19257 1595 19565 1604
rect 2755 1116 3063 1125
rect 2755 1114 2761 1116
rect 2817 1114 2841 1116
rect 2897 1114 2921 1116
rect 2977 1114 3001 1116
rect 3057 1114 3063 1116
rect 2817 1062 2819 1114
rect 2999 1062 3001 1114
rect 2755 1060 2761 1062
rect 2817 1060 2841 1062
rect 2897 1060 2921 1062
rect 2977 1060 3001 1062
rect 3057 1060 3063 1062
rect 2755 1051 3063 1060
rect 7470 1116 7778 1125
rect 7470 1114 7476 1116
rect 7532 1114 7556 1116
rect 7612 1114 7636 1116
rect 7692 1114 7716 1116
rect 7772 1114 7778 1116
rect 7532 1062 7534 1114
rect 7714 1062 7716 1114
rect 7470 1060 7476 1062
rect 7532 1060 7556 1062
rect 7612 1060 7636 1062
rect 7692 1060 7716 1062
rect 7772 1060 7778 1062
rect 7470 1051 7778 1060
rect 12185 1116 12493 1125
rect 12185 1114 12191 1116
rect 12247 1114 12271 1116
rect 12327 1114 12351 1116
rect 12407 1114 12431 1116
rect 12487 1114 12493 1116
rect 12247 1062 12249 1114
rect 12429 1062 12431 1114
rect 12185 1060 12191 1062
rect 12247 1060 12271 1062
rect 12327 1060 12351 1062
rect 12407 1060 12431 1062
rect 12487 1060 12493 1062
rect 12185 1051 12493 1060
rect 16900 1116 17208 1125
rect 16900 1114 16906 1116
rect 16962 1114 16986 1116
rect 17042 1114 17066 1116
rect 17122 1114 17146 1116
rect 17202 1114 17208 1116
rect 16962 1062 16964 1114
rect 17144 1062 17146 1114
rect 16900 1060 16906 1062
rect 16962 1060 16986 1062
rect 17042 1060 17066 1062
rect 17122 1060 17146 1062
rect 17202 1060 17208 1062
rect 16900 1051 17208 1060
rect 3792 808 3844 814
rect 3792 750 3844 756
rect 6276 808 6328 814
rect 6276 750 6328 756
rect 8760 808 8812 814
rect 8760 750 8812 756
rect 11244 808 11296 814
rect 11244 750 11296 756
rect 13728 808 13780 814
rect 13728 750 13780 756
rect 16212 808 16264 814
rect 16212 750 16264 756
rect 18696 808 18748 814
rect 18696 750 18748 756
rect 3804 490 3832 750
rect 5112 572 5420 581
rect 5112 570 5118 572
rect 5174 570 5198 572
rect 5254 570 5278 572
rect 5334 570 5358 572
rect 5414 570 5420 572
rect 5174 518 5176 570
rect 5356 518 5358 570
rect 5112 516 5118 518
rect 5174 516 5198 518
rect 5254 516 5278 518
rect 5334 516 5358 518
rect 5414 516 5420 518
rect 5112 507 5420 516
rect 6288 490 6316 750
rect 8772 490 8800 750
rect 9827 572 10135 581
rect 9827 570 9833 572
rect 9889 570 9913 572
rect 9969 570 9993 572
rect 10049 570 10073 572
rect 10129 570 10135 572
rect 9889 518 9891 570
rect 10071 518 10073 570
rect 9827 516 9833 518
rect 9889 516 9913 518
rect 9969 516 9993 518
rect 10049 516 10073 518
rect 10129 516 10135 518
rect 9827 507 10135 516
rect 11256 490 11284 750
rect 13740 490 13768 750
rect 14542 572 14850 581
rect 14542 570 14548 572
rect 14604 570 14628 572
rect 14684 570 14708 572
rect 14764 570 14788 572
rect 14844 570 14850 572
rect 14604 518 14606 570
rect 14786 518 14788 570
rect 14542 516 14548 518
rect 14604 516 14628 518
rect 14684 516 14708 518
rect 14764 516 14788 518
rect 14844 516 14850 518
rect 14542 507 14850 516
rect 16224 490 16252 750
rect 18708 490 18736 750
rect 19257 572 19565 581
rect 19257 570 19263 572
rect 19319 570 19343 572
rect 19399 570 19423 572
rect 19479 570 19503 572
rect 19559 570 19565 572
rect 19319 518 19321 570
rect 19501 518 19503 570
rect 19257 516 19263 518
rect 19319 516 19343 518
rect 19399 516 19423 518
rect 19479 516 19503 518
rect 19559 516 19565 518
rect 19257 507 19565 516
rect 3712 462 3832 490
rect 6196 462 6316 490
rect 8680 462 8800 490
rect 11164 462 11284 490
rect 13648 462 13768 490
rect 16132 462 16252 490
rect 18616 462 18736 490
rect 3712 400 3740 462
rect 6196 400 6224 462
rect 8680 400 8708 462
rect 11164 400 11192 462
rect 13648 400 13676 462
rect 16132 400 16160 462
rect 18616 400 18644 462
rect 1214 0 1270 400
rect 3698 0 3754 400
rect 6182 0 6238 400
rect 8666 0 8722 400
rect 11150 0 11206 400
rect 13634 0 13690 400
rect 16118 0 16174 400
rect 18602 0 18658 400
<< via2 >>
rect 5118 19066 5174 19068
rect 5198 19066 5254 19068
rect 5278 19066 5334 19068
rect 5358 19066 5414 19068
rect 5118 19014 5164 19066
rect 5164 19014 5174 19066
rect 5198 19014 5228 19066
rect 5228 19014 5240 19066
rect 5240 19014 5254 19066
rect 5278 19014 5292 19066
rect 5292 19014 5304 19066
rect 5304 19014 5334 19066
rect 5358 19014 5368 19066
rect 5368 19014 5414 19066
rect 5118 19012 5174 19014
rect 5198 19012 5254 19014
rect 5278 19012 5334 19014
rect 5358 19012 5414 19014
rect 9833 19066 9889 19068
rect 9913 19066 9969 19068
rect 9993 19066 10049 19068
rect 10073 19066 10129 19068
rect 9833 19014 9879 19066
rect 9879 19014 9889 19066
rect 9913 19014 9943 19066
rect 9943 19014 9955 19066
rect 9955 19014 9969 19066
rect 9993 19014 10007 19066
rect 10007 19014 10019 19066
rect 10019 19014 10049 19066
rect 10073 19014 10083 19066
rect 10083 19014 10129 19066
rect 9833 19012 9889 19014
rect 9913 19012 9969 19014
rect 9993 19012 10049 19014
rect 10073 19012 10129 19014
rect 14548 19066 14604 19068
rect 14628 19066 14684 19068
rect 14708 19066 14764 19068
rect 14788 19066 14844 19068
rect 14548 19014 14594 19066
rect 14594 19014 14604 19066
rect 14628 19014 14658 19066
rect 14658 19014 14670 19066
rect 14670 19014 14684 19066
rect 14708 19014 14722 19066
rect 14722 19014 14734 19066
rect 14734 19014 14764 19066
rect 14788 19014 14798 19066
rect 14798 19014 14844 19066
rect 14548 19012 14604 19014
rect 14628 19012 14684 19014
rect 14708 19012 14764 19014
rect 14788 19012 14844 19014
rect 2761 18522 2817 18524
rect 2841 18522 2897 18524
rect 2921 18522 2977 18524
rect 3001 18522 3057 18524
rect 2761 18470 2807 18522
rect 2807 18470 2817 18522
rect 2841 18470 2871 18522
rect 2871 18470 2883 18522
rect 2883 18470 2897 18522
rect 2921 18470 2935 18522
rect 2935 18470 2947 18522
rect 2947 18470 2977 18522
rect 3001 18470 3011 18522
rect 3011 18470 3057 18522
rect 2761 18468 2817 18470
rect 2841 18468 2897 18470
rect 2921 18468 2977 18470
rect 3001 18468 3057 18470
rect 7476 18522 7532 18524
rect 7556 18522 7612 18524
rect 7636 18522 7692 18524
rect 7716 18522 7772 18524
rect 7476 18470 7522 18522
rect 7522 18470 7532 18522
rect 7556 18470 7586 18522
rect 7586 18470 7598 18522
rect 7598 18470 7612 18522
rect 7636 18470 7650 18522
rect 7650 18470 7662 18522
rect 7662 18470 7692 18522
rect 7716 18470 7726 18522
rect 7726 18470 7772 18522
rect 7476 18468 7532 18470
rect 7556 18468 7612 18470
rect 7636 18468 7692 18470
rect 7716 18468 7772 18470
rect 12191 18522 12247 18524
rect 12271 18522 12327 18524
rect 12351 18522 12407 18524
rect 12431 18522 12487 18524
rect 12191 18470 12237 18522
rect 12237 18470 12247 18522
rect 12271 18470 12301 18522
rect 12301 18470 12313 18522
rect 12313 18470 12327 18522
rect 12351 18470 12365 18522
rect 12365 18470 12377 18522
rect 12377 18470 12407 18522
rect 12431 18470 12441 18522
rect 12441 18470 12487 18522
rect 12191 18468 12247 18470
rect 12271 18468 12327 18470
rect 12351 18468 12407 18470
rect 12431 18468 12487 18470
rect 16906 18522 16962 18524
rect 16986 18522 17042 18524
rect 17066 18522 17122 18524
rect 17146 18522 17202 18524
rect 16906 18470 16952 18522
rect 16952 18470 16962 18522
rect 16986 18470 17016 18522
rect 17016 18470 17028 18522
rect 17028 18470 17042 18522
rect 17066 18470 17080 18522
rect 17080 18470 17092 18522
rect 17092 18470 17122 18522
rect 17146 18470 17156 18522
rect 17156 18470 17202 18522
rect 16906 18468 16962 18470
rect 16986 18468 17042 18470
rect 17066 18468 17122 18470
rect 17146 18468 17202 18470
rect 5118 17978 5174 17980
rect 5198 17978 5254 17980
rect 5278 17978 5334 17980
rect 5358 17978 5414 17980
rect 5118 17926 5164 17978
rect 5164 17926 5174 17978
rect 5198 17926 5228 17978
rect 5228 17926 5240 17978
rect 5240 17926 5254 17978
rect 5278 17926 5292 17978
rect 5292 17926 5304 17978
rect 5304 17926 5334 17978
rect 5358 17926 5368 17978
rect 5368 17926 5414 17978
rect 5118 17924 5174 17926
rect 5198 17924 5254 17926
rect 5278 17924 5334 17926
rect 5358 17924 5414 17926
rect 9833 17978 9889 17980
rect 9913 17978 9969 17980
rect 9993 17978 10049 17980
rect 10073 17978 10129 17980
rect 9833 17926 9879 17978
rect 9879 17926 9889 17978
rect 9913 17926 9943 17978
rect 9943 17926 9955 17978
rect 9955 17926 9969 17978
rect 9993 17926 10007 17978
rect 10007 17926 10019 17978
rect 10019 17926 10049 17978
rect 10073 17926 10083 17978
rect 10083 17926 10129 17978
rect 9833 17924 9889 17926
rect 9913 17924 9969 17926
rect 9993 17924 10049 17926
rect 10073 17924 10129 17926
rect 2761 17434 2817 17436
rect 2841 17434 2897 17436
rect 2921 17434 2977 17436
rect 3001 17434 3057 17436
rect 2761 17382 2807 17434
rect 2807 17382 2817 17434
rect 2841 17382 2871 17434
rect 2871 17382 2883 17434
rect 2883 17382 2897 17434
rect 2921 17382 2935 17434
rect 2935 17382 2947 17434
rect 2947 17382 2977 17434
rect 3001 17382 3011 17434
rect 3011 17382 3057 17434
rect 2761 17380 2817 17382
rect 2841 17380 2897 17382
rect 2921 17380 2977 17382
rect 3001 17380 3057 17382
rect 7476 17434 7532 17436
rect 7556 17434 7612 17436
rect 7636 17434 7692 17436
rect 7716 17434 7772 17436
rect 7476 17382 7522 17434
rect 7522 17382 7532 17434
rect 7556 17382 7586 17434
rect 7586 17382 7598 17434
rect 7598 17382 7612 17434
rect 7636 17382 7650 17434
rect 7650 17382 7662 17434
rect 7662 17382 7692 17434
rect 7716 17382 7726 17434
rect 7726 17382 7772 17434
rect 7476 17380 7532 17382
rect 7556 17380 7612 17382
rect 7636 17380 7692 17382
rect 7716 17380 7772 17382
rect 12191 17434 12247 17436
rect 12271 17434 12327 17436
rect 12351 17434 12407 17436
rect 12431 17434 12487 17436
rect 12191 17382 12237 17434
rect 12237 17382 12247 17434
rect 12271 17382 12301 17434
rect 12301 17382 12313 17434
rect 12313 17382 12327 17434
rect 12351 17382 12365 17434
rect 12365 17382 12377 17434
rect 12377 17382 12407 17434
rect 12431 17382 12441 17434
rect 12441 17382 12487 17434
rect 12191 17380 12247 17382
rect 12271 17380 12327 17382
rect 12351 17380 12407 17382
rect 12431 17380 12487 17382
rect 5118 16890 5174 16892
rect 5198 16890 5254 16892
rect 5278 16890 5334 16892
rect 5358 16890 5414 16892
rect 5118 16838 5164 16890
rect 5164 16838 5174 16890
rect 5198 16838 5228 16890
rect 5228 16838 5240 16890
rect 5240 16838 5254 16890
rect 5278 16838 5292 16890
rect 5292 16838 5304 16890
rect 5304 16838 5334 16890
rect 5358 16838 5368 16890
rect 5368 16838 5414 16890
rect 5118 16836 5174 16838
rect 5198 16836 5254 16838
rect 5278 16836 5334 16838
rect 5358 16836 5414 16838
rect 9833 16890 9889 16892
rect 9913 16890 9969 16892
rect 9993 16890 10049 16892
rect 10073 16890 10129 16892
rect 9833 16838 9879 16890
rect 9879 16838 9889 16890
rect 9913 16838 9943 16890
rect 9943 16838 9955 16890
rect 9955 16838 9969 16890
rect 9993 16838 10007 16890
rect 10007 16838 10019 16890
rect 10019 16838 10049 16890
rect 10073 16838 10083 16890
rect 10083 16838 10129 16890
rect 9833 16836 9889 16838
rect 9913 16836 9969 16838
rect 9993 16836 10049 16838
rect 10073 16836 10129 16838
rect 14548 17978 14604 17980
rect 14628 17978 14684 17980
rect 14708 17978 14764 17980
rect 14788 17978 14844 17980
rect 14548 17926 14594 17978
rect 14594 17926 14604 17978
rect 14628 17926 14658 17978
rect 14658 17926 14670 17978
rect 14670 17926 14684 17978
rect 14708 17926 14722 17978
rect 14722 17926 14734 17978
rect 14734 17926 14764 17978
rect 14788 17926 14798 17978
rect 14798 17926 14844 17978
rect 14548 17924 14604 17926
rect 14628 17924 14684 17926
rect 14708 17924 14764 17926
rect 14788 17924 14844 17926
rect 16906 17434 16962 17436
rect 16986 17434 17042 17436
rect 17066 17434 17122 17436
rect 17146 17434 17202 17436
rect 16906 17382 16952 17434
rect 16952 17382 16962 17434
rect 16986 17382 17016 17434
rect 17016 17382 17028 17434
rect 17028 17382 17042 17434
rect 17066 17382 17080 17434
rect 17080 17382 17092 17434
rect 17092 17382 17122 17434
rect 17146 17382 17156 17434
rect 17156 17382 17202 17434
rect 16906 17380 16962 17382
rect 16986 17380 17042 17382
rect 17066 17380 17122 17382
rect 17146 17380 17202 17382
rect 19263 19066 19319 19068
rect 19343 19066 19399 19068
rect 19423 19066 19479 19068
rect 19503 19066 19559 19068
rect 19263 19014 19309 19066
rect 19309 19014 19319 19066
rect 19343 19014 19373 19066
rect 19373 19014 19385 19066
rect 19385 19014 19399 19066
rect 19423 19014 19437 19066
rect 19437 19014 19449 19066
rect 19449 19014 19479 19066
rect 19503 19014 19513 19066
rect 19513 19014 19559 19066
rect 19263 19012 19319 19014
rect 19343 19012 19399 19014
rect 19423 19012 19479 19014
rect 19503 19012 19559 19014
rect 19263 17978 19319 17980
rect 19343 17978 19399 17980
rect 19423 17978 19479 17980
rect 19503 17978 19559 17980
rect 19263 17926 19309 17978
rect 19309 17926 19319 17978
rect 19343 17926 19373 17978
rect 19373 17926 19385 17978
rect 19385 17926 19399 17978
rect 19423 17926 19437 17978
rect 19437 17926 19449 17978
rect 19449 17926 19479 17978
rect 19503 17926 19513 17978
rect 19513 17926 19559 17978
rect 19263 17924 19319 17926
rect 19343 17924 19399 17926
rect 19423 17924 19479 17926
rect 19503 17924 19559 17926
rect 14548 16890 14604 16892
rect 14628 16890 14684 16892
rect 14708 16890 14764 16892
rect 14788 16890 14844 16892
rect 14548 16838 14594 16890
rect 14594 16838 14604 16890
rect 14628 16838 14658 16890
rect 14658 16838 14670 16890
rect 14670 16838 14684 16890
rect 14708 16838 14722 16890
rect 14722 16838 14734 16890
rect 14734 16838 14764 16890
rect 14788 16838 14798 16890
rect 14798 16838 14844 16890
rect 14548 16836 14604 16838
rect 14628 16836 14684 16838
rect 14708 16836 14764 16838
rect 14788 16836 14844 16838
rect 19263 16890 19319 16892
rect 19343 16890 19399 16892
rect 19423 16890 19479 16892
rect 19503 16890 19559 16892
rect 19263 16838 19309 16890
rect 19309 16838 19319 16890
rect 19343 16838 19373 16890
rect 19373 16838 19385 16890
rect 19385 16838 19399 16890
rect 19423 16838 19437 16890
rect 19437 16838 19449 16890
rect 19449 16838 19479 16890
rect 19503 16838 19513 16890
rect 19513 16838 19559 16890
rect 19263 16836 19319 16838
rect 19343 16836 19399 16838
rect 19423 16836 19479 16838
rect 19503 16836 19559 16838
rect 2761 16346 2817 16348
rect 2841 16346 2897 16348
rect 2921 16346 2977 16348
rect 3001 16346 3057 16348
rect 2761 16294 2807 16346
rect 2807 16294 2817 16346
rect 2841 16294 2871 16346
rect 2871 16294 2883 16346
rect 2883 16294 2897 16346
rect 2921 16294 2935 16346
rect 2935 16294 2947 16346
rect 2947 16294 2977 16346
rect 3001 16294 3011 16346
rect 3011 16294 3057 16346
rect 2761 16292 2817 16294
rect 2841 16292 2897 16294
rect 2921 16292 2977 16294
rect 3001 16292 3057 16294
rect 7476 16346 7532 16348
rect 7556 16346 7612 16348
rect 7636 16346 7692 16348
rect 7716 16346 7772 16348
rect 7476 16294 7522 16346
rect 7522 16294 7532 16346
rect 7556 16294 7586 16346
rect 7586 16294 7598 16346
rect 7598 16294 7612 16346
rect 7636 16294 7650 16346
rect 7650 16294 7662 16346
rect 7662 16294 7692 16346
rect 7716 16294 7726 16346
rect 7726 16294 7772 16346
rect 7476 16292 7532 16294
rect 7556 16292 7612 16294
rect 7636 16292 7692 16294
rect 7716 16292 7772 16294
rect 12191 16346 12247 16348
rect 12271 16346 12327 16348
rect 12351 16346 12407 16348
rect 12431 16346 12487 16348
rect 12191 16294 12237 16346
rect 12237 16294 12247 16346
rect 12271 16294 12301 16346
rect 12301 16294 12313 16346
rect 12313 16294 12327 16346
rect 12351 16294 12365 16346
rect 12365 16294 12377 16346
rect 12377 16294 12407 16346
rect 12431 16294 12441 16346
rect 12441 16294 12487 16346
rect 12191 16292 12247 16294
rect 12271 16292 12327 16294
rect 12351 16292 12407 16294
rect 12431 16292 12487 16294
rect 16906 16346 16962 16348
rect 16986 16346 17042 16348
rect 17066 16346 17122 16348
rect 17146 16346 17202 16348
rect 16906 16294 16952 16346
rect 16952 16294 16962 16346
rect 16986 16294 17016 16346
rect 17016 16294 17028 16346
rect 17028 16294 17042 16346
rect 17066 16294 17080 16346
rect 17080 16294 17092 16346
rect 17092 16294 17122 16346
rect 17146 16294 17156 16346
rect 17156 16294 17202 16346
rect 16906 16292 16962 16294
rect 16986 16292 17042 16294
rect 17066 16292 17122 16294
rect 17146 16292 17202 16294
rect 5118 15802 5174 15804
rect 5198 15802 5254 15804
rect 5278 15802 5334 15804
rect 5358 15802 5414 15804
rect 5118 15750 5164 15802
rect 5164 15750 5174 15802
rect 5198 15750 5228 15802
rect 5228 15750 5240 15802
rect 5240 15750 5254 15802
rect 5278 15750 5292 15802
rect 5292 15750 5304 15802
rect 5304 15750 5334 15802
rect 5358 15750 5368 15802
rect 5368 15750 5414 15802
rect 5118 15748 5174 15750
rect 5198 15748 5254 15750
rect 5278 15748 5334 15750
rect 5358 15748 5414 15750
rect 9833 15802 9889 15804
rect 9913 15802 9969 15804
rect 9993 15802 10049 15804
rect 10073 15802 10129 15804
rect 9833 15750 9879 15802
rect 9879 15750 9889 15802
rect 9913 15750 9943 15802
rect 9943 15750 9955 15802
rect 9955 15750 9969 15802
rect 9993 15750 10007 15802
rect 10007 15750 10019 15802
rect 10019 15750 10049 15802
rect 10073 15750 10083 15802
rect 10083 15750 10129 15802
rect 9833 15748 9889 15750
rect 9913 15748 9969 15750
rect 9993 15748 10049 15750
rect 10073 15748 10129 15750
rect 14548 15802 14604 15804
rect 14628 15802 14684 15804
rect 14708 15802 14764 15804
rect 14788 15802 14844 15804
rect 14548 15750 14594 15802
rect 14594 15750 14604 15802
rect 14628 15750 14658 15802
rect 14658 15750 14670 15802
rect 14670 15750 14684 15802
rect 14708 15750 14722 15802
rect 14722 15750 14734 15802
rect 14734 15750 14764 15802
rect 14788 15750 14798 15802
rect 14798 15750 14844 15802
rect 14548 15748 14604 15750
rect 14628 15748 14684 15750
rect 14708 15748 14764 15750
rect 14788 15748 14844 15750
rect 19263 15802 19319 15804
rect 19343 15802 19399 15804
rect 19423 15802 19479 15804
rect 19503 15802 19559 15804
rect 19263 15750 19309 15802
rect 19309 15750 19319 15802
rect 19343 15750 19373 15802
rect 19373 15750 19385 15802
rect 19385 15750 19399 15802
rect 19423 15750 19437 15802
rect 19437 15750 19449 15802
rect 19449 15750 19479 15802
rect 19503 15750 19513 15802
rect 19513 15750 19559 15802
rect 19263 15748 19319 15750
rect 19343 15748 19399 15750
rect 19423 15748 19479 15750
rect 19503 15748 19559 15750
rect 2761 15258 2817 15260
rect 2841 15258 2897 15260
rect 2921 15258 2977 15260
rect 3001 15258 3057 15260
rect 2761 15206 2807 15258
rect 2807 15206 2817 15258
rect 2841 15206 2871 15258
rect 2871 15206 2883 15258
rect 2883 15206 2897 15258
rect 2921 15206 2935 15258
rect 2935 15206 2947 15258
rect 2947 15206 2977 15258
rect 3001 15206 3011 15258
rect 3011 15206 3057 15258
rect 2761 15204 2817 15206
rect 2841 15204 2897 15206
rect 2921 15204 2977 15206
rect 3001 15204 3057 15206
rect 7476 15258 7532 15260
rect 7556 15258 7612 15260
rect 7636 15258 7692 15260
rect 7716 15258 7772 15260
rect 7476 15206 7522 15258
rect 7522 15206 7532 15258
rect 7556 15206 7586 15258
rect 7586 15206 7598 15258
rect 7598 15206 7612 15258
rect 7636 15206 7650 15258
rect 7650 15206 7662 15258
rect 7662 15206 7692 15258
rect 7716 15206 7726 15258
rect 7726 15206 7772 15258
rect 7476 15204 7532 15206
rect 7556 15204 7612 15206
rect 7636 15204 7692 15206
rect 7716 15204 7772 15206
rect 12191 15258 12247 15260
rect 12271 15258 12327 15260
rect 12351 15258 12407 15260
rect 12431 15258 12487 15260
rect 12191 15206 12237 15258
rect 12237 15206 12247 15258
rect 12271 15206 12301 15258
rect 12301 15206 12313 15258
rect 12313 15206 12327 15258
rect 12351 15206 12365 15258
rect 12365 15206 12377 15258
rect 12377 15206 12407 15258
rect 12431 15206 12441 15258
rect 12441 15206 12487 15258
rect 12191 15204 12247 15206
rect 12271 15204 12327 15206
rect 12351 15204 12407 15206
rect 12431 15204 12487 15206
rect 16906 15258 16962 15260
rect 16986 15258 17042 15260
rect 17066 15258 17122 15260
rect 17146 15258 17202 15260
rect 16906 15206 16952 15258
rect 16952 15206 16962 15258
rect 16986 15206 17016 15258
rect 17016 15206 17028 15258
rect 17028 15206 17042 15258
rect 17066 15206 17080 15258
rect 17080 15206 17092 15258
rect 17092 15206 17122 15258
rect 17146 15206 17156 15258
rect 17156 15206 17202 15258
rect 16906 15204 16962 15206
rect 16986 15204 17042 15206
rect 17066 15204 17122 15206
rect 17146 15204 17202 15206
rect 5118 14714 5174 14716
rect 5198 14714 5254 14716
rect 5278 14714 5334 14716
rect 5358 14714 5414 14716
rect 5118 14662 5164 14714
rect 5164 14662 5174 14714
rect 5198 14662 5228 14714
rect 5228 14662 5240 14714
rect 5240 14662 5254 14714
rect 5278 14662 5292 14714
rect 5292 14662 5304 14714
rect 5304 14662 5334 14714
rect 5358 14662 5368 14714
rect 5368 14662 5414 14714
rect 5118 14660 5174 14662
rect 5198 14660 5254 14662
rect 5278 14660 5334 14662
rect 5358 14660 5414 14662
rect 9833 14714 9889 14716
rect 9913 14714 9969 14716
rect 9993 14714 10049 14716
rect 10073 14714 10129 14716
rect 9833 14662 9879 14714
rect 9879 14662 9889 14714
rect 9913 14662 9943 14714
rect 9943 14662 9955 14714
rect 9955 14662 9969 14714
rect 9993 14662 10007 14714
rect 10007 14662 10019 14714
rect 10019 14662 10049 14714
rect 10073 14662 10083 14714
rect 10083 14662 10129 14714
rect 9833 14660 9889 14662
rect 9913 14660 9969 14662
rect 9993 14660 10049 14662
rect 10073 14660 10129 14662
rect 14548 14714 14604 14716
rect 14628 14714 14684 14716
rect 14708 14714 14764 14716
rect 14788 14714 14844 14716
rect 14548 14662 14594 14714
rect 14594 14662 14604 14714
rect 14628 14662 14658 14714
rect 14658 14662 14670 14714
rect 14670 14662 14684 14714
rect 14708 14662 14722 14714
rect 14722 14662 14734 14714
rect 14734 14662 14764 14714
rect 14788 14662 14798 14714
rect 14798 14662 14844 14714
rect 14548 14660 14604 14662
rect 14628 14660 14684 14662
rect 14708 14660 14764 14662
rect 14788 14660 14844 14662
rect 19263 14714 19319 14716
rect 19343 14714 19399 14716
rect 19423 14714 19479 14716
rect 19503 14714 19559 14716
rect 19263 14662 19309 14714
rect 19309 14662 19319 14714
rect 19343 14662 19373 14714
rect 19373 14662 19385 14714
rect 19385 14662 19399 14714
rect 19423 14662 19437 14714
rect 19437 14662 19449 14714
rect 19449 14662 19479 14714
rect 19503 14662 19513 14714
rect 19513 14662 19559 14714
rect 19263 14660 19319 14662
rect 19343 14660 19399 14662
rect 19423 14660 19479 14662
rect 19503 14660 19559 14662
rect 2761 14170 2817 14172
rect 2841 14170 2897 14172
rect 2921 14170 2977 14172
rect 3001 14170 3057 14172
rect 2761 14118 2807 14170
rect 2807 14118 2817 14170
rect 2841 14118 2871 14170
rect 2871 14118 2883 14170
rect 2883 14118 2897 14170
rect 2921 14118 2935 14170
rect 2935 14118 2947 14170
rect 2947 14118 2977 14170
rect 3001 14118 3011 14170
rect 3011 14118 3057 14170
rect 2761 14116 2817 14118
rect 2841 14116 2897 14118
rect 2921 14116 2977 14118
rect 3001 14116 3057 14118
rect 7476 14170 7532 14172
rect 7556 14170 7612 14172
rect 7636 14170 7692 14172
rect 7716 14170 7772 14172
rect 7476 14118 7522 14170
rect 7522 14118 7532 14170
rect 7556 14118 7586 14170
rect 7586 14118 7598 14170
rect 7598 14118 7612 14170
rect 7636 14118 7650 14170
rect 7650 14118 7662 14170
rect 7662 14118 7692 14170
rect 7716 14118 7726 14170
rect 7726 14118 7772 14170
rect 7476 14116 7532 14118
rect 7556 14116 7612 14118
rect 7636 14116 7692 14118
rect 7716 14116 7772 14118
rect 12191 14170 12247 14172
rect 12271 14170 12327 14172
rect 12351 14170 12407 14172
rect 12431 14170 12487 14172
rect 12191 14118 12237 14170
rect 12237 14118 12247 14170
rect 12271 14118 12301 14170
rect 12301 14118 12313 14170
rect 12313 14118 12327 14170
rect 12351 14118 12365 14170
rect 12365 14118 12377 14170
rect 12377 14118 12407 14170
rect 12431 14118 12441 14170
rect 12441 14118 12487 14170
rect 12191 14116 12247 14118
rect 12271 14116 12327 14118
rect 12351 14116 12407 14118
rect 12431 14116 12487 14118
rect 16906 14170 16962 14172
rect 16986 14170 17042 14172
rect 17066 14170 17122 14172
rect 17146 14170 17202 14172
rect 16906 14118 16952 14170
rect 16952 14118 16962 14170
rect 16986 14118 17016 14170
rect 17016 14118 17028 14170
rect 17028 14118 17042 14170
rect 17066 14118 17080 14170
rect 17080 14118 17092 14170
rect 17092 14118 17122 14170
rect 17146 14118 17156 14170
rect 17156 14118 17202 14170
rect 16906 14116 16962 14118
rect 16986 14116 17042 14118
rect 17066 14116 17122 14118
rect 17146 14116 17202 14118
rect 5118 13626 5174 13628
rect 5198 13626 5254 13628
rect 5278 13626 5334 13628
rect 5358 13626 5414 13628
rect 5118 13574 5164 13626
rect 5164 13574 5174 13626
rect 5198 13574 5228 13626
rect 5228 13574 5240 13626
rect 5240 13574 5254 13626
rect 5278 13574 5292 13626
rect 5292 13574 5304 13626
rect 5304 13574 5334 13626
rect 5358 13574 5368 13626
rect 5368 13574 5414 13626
rect 5118 13572 5174 13574
rect 5198 13572 5254 13574
rect 5278 13572 5334 13574
rect 5358 13572 5414 13574
rect 9833 13626 9889 13628
rect 9913 13626 9969 13628
rect 9993 13626 10049 13628
rect 10073 13626 10129 13628
rect 9833 13574 9879 13626
rect 9879 13574 9889 13626
rect 9913 13574 9943 13626
rect 9943 13574 9955 13626
rect 9955 13574 9969 13626
rect 9993 13574 10007 13626
rect 10007 13574 10019 13626
rect 10019 13574 10049 13626
rect 10073 13574 10083 13626
rect 10083 13574 10129 13626
rect 9833 13572 9889 13574
rect 9913 13572 9969 13574
rect 9993 13572 10049 13574
rect 10073 13572 10129 13574
rect 14548 13626 14604 13628
rect 14628 13626 14684 13628
rect 14708 13626 14764 13628
rect 14788 13626 14844 13628
rect 14548 13574 14594 13626
rect 14594 13574 14604 13626
rect 14628 13574 14658 13626
rect 14658 13574 14670 13626
rect 14670 13574 14684 13626
rect 14708 13574 14722 13626
rect 14722 13574 14734 13626
rect 14734 13574 14764 13626
rect 14788 13574 14798 13626
rect 14798 13574 14844 13626
rect 14548 13572 14604 13574
rect 14628 13572 14684 13574
rect 14708 13572 14764 13574
rect 14788 13572 14844 13574
rect 19263 13626 19319 13628
rect 19343 13626 19399 13628
rect 19423 13626 19479 13628
rect 19503 13626 19559 13628
rect 19263 13574 19309 13626
rect 19309 13574 19319 13626
rect 19343 13574 19373 13626
rect 19373 13574 19385 13626
rect 19385 13574 19399 13626
rect 19423 13574 19437 13626
rect 19437 13574 19449 13626
rect 19449 13574 19479 13626
rect 19503 13574 19513 13626
rect 19513 13574 19559 13626
rect 19263 13572 19319 13574
rect 19343 13572 19399 13574
rect 19423 13572 19479 13574
rect 19503 13572 19559 13574
rect 2761 13082 2817 13084
rect 2841 13082 2897 13084
rect 2921 13082 2977 13084
rect 3001 13082 3057 13084
rect 2761 13030 2807 13082
rect 2807 13030 2817 13082
rect 2841 13030 2871 13082
rect 2871 13030 2883 13082
rect 2883 13030 2897 13082
rect 2921 13030 2935 13082
rect 2935 13030 2947 13082
rect 2947 13030 2977 13082
rect 3001 13030 3011 13082
rect 3011 13030 3057 13082
rect 2761 13028 2817 13030
rect 2841 13028 2897 13030
rect 2921 13028 2977 13030
rect 3001 13028 3057 13030
rect 7476 13082 7532 13084
rect 7556 13082 7612 13084
rect 7636 13082 7692 13084
rect 7716 13082 7772 13084
rect 7476 13030 7522 13082
rect 7522 13030 7532 13082
rect 7556 13030 7586 13082
rect 7586 13030 7598 13082
rect 7598 13030 7612 13082
rect 7636 13030 7650 13082
rect 7650 13030 7662 13082
rect 7662 13030 7692 13082
rect 7716 13030 7726 13082
rect 7726 13030 7772 13082
rect 7476 13028 7532 13030
rect 7556 13028 7612 13030
rect 7636 13028 7692 13030
rect 7716 13028 7772 13030
rect 12191 13082 12247 13084
rect 12271 13082 12327 13084
rect 12351 13082 12407 13084
rect 12431 13082 12487 13084
rect 12191 13030 12237 13082
rect 12237 13030 12247 13082
rect 12271 13030 12301 13082
rect 12301 13030 12313 13082
rect 12313 13030 12327 13082
rect 12351 13030 12365 13082
rect 12365 13030 12377 13082
rect 12377 13030 12407 13082
rect 12431 13030 12441 13082
rect 12441 13030 12487 13082
rect 12191 13028 12247 13030
rect 12271 13028 12327 13030
rect 12351 13028 12407 13030
rect 12431 13028 12487 13030
rect 16906 13082 16962 13084
rect 16986 13082 17042 13084
rect 17066 13082 17122 13084
rect 17146 13082 17202 13084
rect 16906 13030 16952 13082
rect 16952 13030 16962 13082
rect 16986 13030 17016 13082
rect 17016 13030 17028 13082
rect 17028 13030 17042 13082
rect 17066 13030 17080 13082
rect 17080 13030 17092 13082
rect 17092 13030 17122 13082
rect 17146 13030 17156 13082
rect 17156 13030 17202 13082
rect 16906 13028 16962 13030
rect 16986 13028 17042 13030
rect 17066 13028 17122 13030
rect 17146 13028 17202 13030
rect 5118 12538 5174 12540
rect 5198 12538 5254 12540
rect 5278 12538 5334 12540
rect 5358 12538 5414 12540
rect 5118 12486 5164 12538
rect 5164 12486 5174 12538
rect 5198 12486 5228 12538
rect 5228 12486 5240 12538
rect 5240 12486 5254 12538
rect 5278 12486 5292 12538
rect 5292 12486 5304 12538
rect 5304 12486 5334 12538
rect 5358 12486 5368 12538
rect 5368 12486 5414 12538
rect 5118 12484 5174 12486
rect 5198 12484 5254 12486
rect 5278 12484 5334 12486
rect 5358 12484 5414 12486
rect 9833 12538 9889 12540
rect 9913 12538 9969 12540
rect 9993 12538 10049 12540
rect 10073 12538 10129 12540
rect 9833 12486 9879 12538
rect 9879 12486 9889 12538
rect 9913 12486 9943 12538
rect 9943 12486 9955 12538
rect 9955 12486 9969 12538
rect 9993 12486 10007 12538
rect 10007 12486 10019 12538
rect 10019 12486 10049 12538
rect 10073 12486 10083 12538
rect 10083 12486 10129 12538
rect 9833 12484 9889 12486
rect 9913 12484 9969 12486
rect 9993 12484 10049 12486
rect 10073 12484 10129 12486
rect 14548 12538 14604 12540
rect 14628 12538 14684 12540
rect 14708 12538 14764 12540
rect 14788 12538 14844 12540
rect 14548 12486 14594 12538
rect 14594 12486 14604 12538
rect 14628 12486 14658 12538
rect 14658 12486 14670 12538
rect 14670 12486 14684 12538
rect 14708 12486 14722 12538
rect 14722 12486 14734 12538
rect 14734 12486 14764 12538
rect 14788 12486 14798 12538
rect 14798 12486 14844 12538
rect 14548 12484 14604 12486
rect 14628 12484 14684 12486
rect 14708 12484 14764 12486
rect 14788 12484 14844 12486
rect 19263 12538 19319 12540
rect 19343 12538 19399 12540
rect 19423 12538 19479 12540
rect 19503 12538 19559 12540
rect 19263 12486 19309 12538
rect 19309 12486 19319 12538
rect 19343 12486 19373 12538
rect 19373 12486 19385 12538
rect 19385 12486 19399 12538
rect 19423 12486 19437 12538
rect 19437 12486 19449 12538
rect 19449 12486 19479 12538
rect 19503 12486 19513 12538
rect 19513 12486 19559 12538
rect 19263 12484 19319 12486
rect 19343 12484 19399 12486
rect 19423 12484 19479 12486
rect 19503 12484 19559 12486
rect 2761 11994 2817 11996
rect 2841 11994 2897 11996
rect 2921 11994 2977 11996
rect 3001 11994 3057 11996
rect 2761 11942 2807 11994
rect 2807 11942 2817 11994
rect 2841 11942 2871 11994
rect 2871 11942 2883 11994
rect 2883 11942 2897 11994
rect 2921 11942 2935 11994
rect 2935 11942 2947 11994
rect 2947 11942 2977 11994
rect 3001 11942 3011 11994
rect 3011 11942 3057 11994
rect 2761 11940 2817 11942
rect 2841 11940 2897 11942
rect 2921 11940 2977 11942
rect 3001 11940 3057 11942
rect 7476 11994 7532 11996
rect 7556 11994 7612 11996
rect 7636 11994 7692 11996
rect 7716 11994 7772 11996
rect 7476 11942 7522 11994
rect 7522 11942 7532 11994
rect 7556 11942 7586 11994
rect 7586 11942 7598 11994
rect 7598 11942 7612 11994
rect 7636 11942 7650 11994
rect 7650 11942 7662 11994
rect 7662 11942 7692 11994
rect 7716 11942 7726 11994
rect 7726 11942 7772 11994
rect 7476 11940 7532 11942
rect 7556 11940 7612 11942
rect 7636 11940 7692 11942
rect 7716 11940 7772 11942
rect 12191 11994 12247 11996
rect 12271 11994 12327 11996
rect 12351 11994 12407 11996
rect 12431 11994 12487 11996
rect 12191 11942 12237 11994
rect 12237 11942 12247 11994
rect 12271 11942 12301 11994
rect 12301 11942 12313 11994
rect 12313 11942 12327 11994
rect 12351 11942 12365 11994
rect 12365 11942 12377 11994
rect 12377 11942 12407 11994
rect 12431 11942 12441 11994
rect 12441 11942 12487 11994
rect 12191 11940 12247 11942
rect 12271 11940 12327 11942
rect 12351 11940 12407 11942
rect 12431 11940 12487 11942
rect 16906 11994 16962 11996
rect 16986 11994 17042 11996
rect 17066 11994 17122 11996
rect 17146 11994 17202 11996
rect 16906 11942 16952 11994
rect 16952 11942 16962 11994
rect 16986 11942 17016 11994
rect 17016 11942 17028 11994
rect 17028 11942 17042 11994
rect 17066 11942 17080 11994
rect 17080 11942 17092 11994
rect 17092 11942 17122 11994
rect 17146 11942 17156 11994
rect 17156 11942 17202 11994
rect 16906 11940 16962 11942
rect 16986 11940 17042 11942
rect 17066 11940 17122 11942
rect 17146 11940 17202 11942
rect 5118 11450 5174 11452
rect 5198 11450 5254 11452
rect 5278 11450 5334 11452
rect 5358 11450 5414 11452
rect 5118 11398 5164 11450
rect 5164 11398 5174 11450
rect 5198 11398 5228 11450
rect 5228 11398 5240 11450
rect 5240 11398 5254 11450
rect 5278 11398 5292 11450
rect 5292 11398 5304 11450
rect 5304 11398 5334 11450
rect 5358 11398 5368 11450
rect 5368 11398 5414 11450
rect 5118 11396 5174 11398
rect 5198 11396 5254 11398
rect 5278 11396 5334 11398
rect 5358 11396 5414 11398
rect 9833 11450 9889 11452
rect 9913 11450 9969 11452
rect 9993 11450 10049 11452
rect 10073 11450 10129 11452
rect 9833 11398 9879 11450
rect 9879 11398 9889 11450
rect 9913 11398 9943 11450
rect 9943 11398 9955 11450
rect 9955 11398 9969 11450
rect 9993 11398 10007 11450
rect 10007 11398 10019 11450
rect 10019 11398 10049 11450
rect 10073 11398 10083 11450
rect 10083 11398 10129 11450
rect 9833 11396 9889 11398
rect 9913 11396 9969 11398
rect 9993 11396 10049 11398
rect 10073 11396 10129 11398
rect 14548 11450 14604 11452
rect 14628 11450 14684 11452
rect 14708 11450 14764 11452
rect 14788 11450 14844 11452
rect 14548 11398 14594 11450
rect 14594 11398 14604 11450
rect 14628 11398 14658 11450
rect 14658 11398 14670 11450
rect 14670 11398 14684 11450
rect 14708 11398 14722 11450
rect 14722 11398 14734 11450
rect 14734 11398 14764 11450
rect 14788 11398 14798 11450
rect 14798 11398 14844 11450
rect 14548 11396 14604 11398
rect 14628 11396 14684 11398
rect 14708 11396 14764 11398
rect 14788 11396 14844 11398
rect 19263 11450 19319 11452
rect 19343 11450 19399 11452
rect 19423 11450 19479 11452
rect 19503 11450 19559 11452
rect 19263 11398 19309 11450
rect 19309 11398 19319 11450
rect 19343 11398 19373 11450
rect 19373 11398 19385 11450
rect 19385 11398 19399 11450
rect 19423 11398 19437 11450
rect 19437 11398 19449 11450
rect 19449 11398 19479 11450
rect 19503 11398 19513 11450
rect 19513 11398 19559 11450
rect 19263 11396 19319 11398
rect 19343 11396 19399 11398
rect 19423 11396 19479 11398
rect 19503 11396 19559 11398
rect 2761 10906 2817 10908
rect 2841 10906 2897 10908
rect 2921 10906 2977 10908
rect 3001 10906 3057 10908
rect 2761 10854 2807 10906
rect 2807 10854 2817 10906
rect 2841 10854 2871 10906
rect 2871 10854 2883 10906
rect 2883 10854 2897 10906
rect 2921 10854 2935 10906
rect 2935 10854 2947 10906
rect 2947 10854 2977 10906
rect 3001 10854 3011 10906
rect 3011 10854 3057 10906
rect 2761 10852 2817 10854
rect 2841 10852 2897 10854
rect 2921 10852 2977 10854
rect 3001 10852 3057 10854
rect 7476 10906 7532 10908
rect 7556 10906 7612 10908
rect 7636 10906 7692 10908
rect 7716 10906 7772 10908
rect 7476 10854 7522 10906
rect 7522 10854 7532 10906
rect 7556 10854 7586 10906
rect 7586 10854 7598 10906
rect 7598 10854 7612 10906
rect 7636 10854 7650 10906
rect 7650 10854 7662 10906
rect 7662 10854 7692 10906
rect 7716 10854 7726 10906
rect 7726 10854 7772 10906
rect 7476 10852 7532 10854
rect 7556 10852 7612 10854
rect 7636 10852 7692 10854
rect 7716 10852 7772 10854
rect 12191 10906 12247 10908
rect 12271 10906 12327 10908
rect 12351 10906 12407 10908
rect 12431 10906 12487 10908
rect 12191 10854 12237 10906
rect 12237 10854 12247 10906
rect 12271 10854 12301 10906
rect 12301 10854 12313 10906
rect 12313 10854 12327 10906
rect 12351 10854 12365 10906
rect 12365 10854 12377 10906
rect 12377 10854 12407 10906
rect 12431 10854 12441 10906
rect 12441 10854 12487 10906
rect 12191 10852 12247 10854
rect 12271 10852 12327 10854
rect 12351 10852 12407 10854
rect 12431 10852 12487 10854
rect 16906 10906 16962 10908
rect 16986 10906 17042 10908
rect 17066 10906 17122 10908
rect 17146 10906 17202 10908
rect 16906 10854 16952 10906
rect 16952 10854 16962 10906
rect 16986 10854 17016 10906
rect 17016 10854 17028 10906
rect 17028 10854 17042 10906
rect 17066 10854 17080 10906
rect 17080 10854 17092 10906
rect 17092 10854 17122 10906
rect 17146 10854 17156 10906
rect 17156 10854 17202 10906
rect 16906 10852 16962 10854
rect 16986 10852 17042 10854
rect 17066 10852 17122 10854
rect 17146 10852 17202 10854
rect 5118 10362 5174 10364
rect 5198 10362 5254 10364
rect 5278 10362 5334 10364
rect 5358 10362 5414 10364
rect 5118 10310 5164 10362
rect 5164 10310 5174 10362
rect 5198 10310 5228 10362
rect 5228 10310 5240 10362
rect 5240 10310 5254 10362
rect 5278 10310 5292 10362
rect 5292 10310 5304 10362
rect 5304 10310 5334 10362
rect 5358 10310 5368 10362
rect 5368 10310 5414 10362
rect 5118 10308 5174 10310
rect 5198 10308 5254 10310
rect 5278 10308 5334 10310
rect 5358 10308 5414 10310
rect 9833 10362 9889 10364
rect 9913 10362 9969 10364
rect 9993 10362 10049 10364
rect 10073 10362 10129 10364
rect 9833 10310 9879 10362
rect 9879 10310 9889 10362
rect 9913 10310 9943 10362
rect 9943 10310 9955 10362
rect 9955 10310 9969 10362
rect 9993 10310 10007 10362
rect 10007 10310 10019 10362
rect 10019 10310 10049 10362
rect 10073 10310 10083 10362
rect 10083 10310 10129 10362
rect 9833 10308 9889 10310
rect 9913 10308 9969 10310
rect 9993 10308 10049 10310
rect 10073 10308 10129 10310
rect 14548 10362 14604 10364
rect 14628 10362 14684 10364
rect 14708 10362 14764 10364
rect 14788 10362 14844 10364
rect 14548 10310 14594 10362
rect 14594 10310 14604 10362
rect 14628 10310 14658 10362
rect 14658 10310 14670 10362
rect 14670 10310 14684 10362
rect 14708 10310 14722 10362
rect 14722 10310 14734 10362
rect 14734 10310 14764 10362
rect 14788 10310 14798 10362
rect 14798 10310 14844 10362
rect 14548 10308 14604 10310
rect 14628 10308 14684 10310
rect 14708 10308 14764 10310
rect 14788 10308 14844 10310
rect 19263 10362 19319 10364
rect 19343 10362 19399 10364
rect 19423 10362 19479 10364
rect 19503 10362 19559 10364
rect 19263 10310 19309 10362
rect 19309 10310 19319 10362
rect 19343 10310 19373 10362
rect 19373 10310 19385 10362
rect 19385 10310 19399 10362
rect 19423 10310 19437 10362
rect 19437 10310 19449 10362
rect 19449 10310 19479 10362
rect 19503 10310 19513 10362
rect 19513 10310 19559 10362
rect 19263 10308 19319 10310
rect 19343 10308 19399 10310
rect 19423 10308 19479 10310
rect 19503 10308 19559 10310
rect 19062 9868 19064 9888
rect 19064 9868 19116 9888
rect 19116 9868 19118 9888
rect 19062 9832 19118 9868
rect 2761 9818 2817 9820
rect 2841 9818 2897 9820
rect 2921 9818 2977 9820
rect 3001 9818 3057 9820
rect 2761 9766 2807 9818
rect 2807 9766 2817 9818
rect 2841 9766 2871 9818
rect 2871 9766 2883 9818
rect 2883 9766 2897 9818
rect 2921 9766 2935 9818
rect 2935 9766 2947 9818
rect 2947 9766 2977 9818
rect 3001 9766 3011 9818
rect 3011 9766 3057 9818
rect 2761 9764 2817 9766
rect 2841 9764 2897 9766
rect 2921 9764 2977 9766
rect 3001 9764 3057 9766
rect 7476 9818 7532 9820
rect 7556 9818 7612 9820
rect 7636 9818 7692 9820
rect 7716 9818 7772 9820
rect 7476 9766 7522 9818
rect 7522 9766 7532 9818
rect 7556 9766 7586 9818
rect 7586 9766 7598 9818
rect 7598 9766 7612 9818
rect 7636 9766 7650 9818
rect 7650 9766 7662 9818
rect 7662 9766 7692 9818
rect 7716 9766 7726 9818
rect 7726 9766 7772 9818
rect 7476 9764 7532 9766
rect 7556 9764 7612 9766
rect 7636 9764 7692 9766
rect 7716 9764 7772 9766
rect 12191 9818 12247 9820
rect 12271 9818 12327 9820
rect 12351 9818 12407 9820
rect 12431 9818 12487 9820
rect 12191 9766 12237 9818
rect 12237 9766 12247 9818
rect 12271 9766 12301 9818
rect 12301 9766 12313 9818
rect 12313 9766 12327 9818
rect 12351 9766 12365 9818
rect 12365 9766 12377 9818
rect 12377 9766 12407 9818
rect 12431 9766 12441 9818
rect 12441 9766 12487 9818
rect 12191 9764 12247 9766
rect 12271 9764 12327 9766
rect 12351 9764 12407 9766
rect 12431 9764 12487 9766
rect 16906 9818 16962 9820
rect 16986 9818 17042 9820
rect 17066 9818 17122 9820
rect 17146 9818 17202 9820
rect 16906 9766 16952 9818
rect 16952 9766 16962 9818
rect 16986 9766 17016 9818
rect 17016 9766 17028 9818
rect 17028 9766 17042 9818
rect 17066 9766 17080 9818
rect 17080 9766 17092 9818
rect 17092 9766 17122 9818
rect 17146 9766 17156 9818
rect 17156 9766 17202 9818
rect 16906 9764 16962 9766
rect 16986 9764 17042 9766
rect 17066 9764 17122 9766
rect 17146 9764 17202 9766
rect 5118 9274 5174 9276
rect 5198 9274 5254 9276
rect 5278 9274 5334 9276
rect 5358 9274 5414 9276
rect 5118 9222 5164 9274
rect 5164 9222 5174 9274
rect 5198 9222 5228 9274
rect 5228 9222 5240 9274
rect 5240 9222 5254 9274
rect 5278 9222 5292 9274
rect 5292 9222 5304 9274
rect 5304 9222 5334 9274
rect 5358 9222 5368 9274
rect 5368 9222 5414 9274
rect 5118 9220 5174 9222
rect 5198 9220 5254 9222
rect 5278 9220 5334 9222
rect 5358 9220 5414 9222
rect 9833 9274 9889 9276
rect 9913 9274 9969 9276
rect 9993 9274 10049 9276
rect 10073 9274 10129 9276
rect 9833 9222 9879 9274
rect 9879 9222 9889 9274
rect 9913 9222 9943 9274
rect 9943 9222 9955 9274
rect 9955 9222 9969 9274
rect 9993 9222 10007 9274
rect 10007 9222 10019 9274
rect 10019 9222 10049 9274
rect 10073 9222 10083 9274
rect 10083 9222 10129 9274
rect 9833 9220 9889 9222
rect 9913 9220 9969 9222
rect 9993 9220 10049 9222
rect 10073 9220 10129 9222
rect 14548 9274 14604 9276
rect 14628 9274 14684 9276
rect 14708 9274 14764 9276
rect 14788 9274 14844 9276
rect 14548 9222 14594 9274
rect 14594 9222 14604 9274
rect 14628 9222 14658 9274
rect 14658 9222 14670 9274
rect 14670 9222 14684 9274
rect 14708 9222 14722 9274
rect 14722 9222 14734 9274
rect 14734 9222 14764 9274
rect 14788 9222 14798 9274
rect 14798 9222 14844 9274
rect 14548 9220 14604 9222
rect 14628 9220 14684 9222
rect 14708 9220 14764 9222
rect 14788 9220 14844 9222
rect 19263 9274 19319 9276
rect 19343 9274 19399 9276
rect 19423 9274 19479 9276
rect 19503 9274 19559 9276
rect 19263 9222 19309 9274
rect 19309 9222 19319 9274
rect 19343 9222 19373 9274
rect 19373 9222 19385 9274
rect 19385 9222 19399 9274
rect 19423 9222 19437 9274
rect 19437 9222 19449 9274
rect 19449 9222 19479 9274
rect 19503 9222 19513 9274
rect 19513 9222 19559 9274
rect 19263 9220 19319 9222
rect 19343 9220 19399 9222
rect 19423 9220 19479 9222
rect 19503 9220 19559 9222
rect 2761 8730 2817 8732
rect 2841 8730 2897 8732
rect 2921 8730 2977 8732
rect 3001 8730 3057 8732
rect 2761 8678 2807 8730
rect 2807 8678 2817 8730
rect 2841 8678 2871 8730
rect 2871 8678 2883 8730
rect 2883 8678 2897 8730
rect 2921 8678 2935 8730
rect 2935 8678 2947 8730
rect 2947 8678 2977 8730
rect 3001 8678 3011 8730
rect 3011 8678 3057 8730
rect 2761 8676 2817 8678
rect 2841 8676 2897 8678
rect 2921 8676 2977 8678
rect 3001 8676 3057 8678
rect 7476 8730 7532 8732
rect 7556 8730 7612 8732
rect 7636 8730 7692 8732
rect 7716 8730 7772 8732
rect 7476 8678 7522 8730
rect 7522 8678 7532 8730
rect 7556 8678 7586 8730
rect 7586 8678 7598 8730
rect 7598 8678 7612 8730
rect 7636 8678 7650 8730
rect 7650 8678 7662 8730
rect 7662 8678 7692 8730
rect 7716 8678 7726 8730
rect 7726 8678 7772 8730
rect 7476 8676 7532 8678
rect 7556 8676 7612 8678
rect 7636 8676 7692 8678
rect 7716 8676 7772 8678
rect 12191 8730 12247 8732
rect 12271 8730 12327 8732
rect 12351 8730 12407 8732
rect 12431 8730 12487 8732
rect 12191 8678 12237 8730
rect 12237 8678 12247 8730
rect 12271 8678 12301 8730
rect 12301 8678 12313 8730
rect 12313 8678 12327 8730
rect 12351 8678 12365 8730
rect 12365 8678 12377 8730
rect 12377 8678 12407 8730
rect 12431 8678 12441 8730
rect 12441 8678 12487 8730
rect 12191 8676 12247 8678
rect 12271 8676 12327 8678
rect 12351 8676 12407 8678
rect 12431 8676 12487 8678
rect 16906 8730 16962 8732
rect 16986 8730 17042 8732
rect 17066 8730 17122 8732
rect 17146 8730 17202 8732
rect 16906 8678 16952 8730
rect 16952 8678 16962 8730
rect 16986 8678 17016 8730
rect 17016 8678 17028 8730
rect 17028 8678 17042 8730
rect 17066 8678 17080 8730
rect 17080 8678 17092 8730
rect 17092 8678 17122 8730
rect 17146 8678 17156 8730
rect 17156 8678 17202 8730
rect 16906 8676 16962 8678
rect 16986 8676 17042 8678
rect 17066 8676 17122 8678
rect 17146 8676 17202 8678
rect 5118 8186 5174 8188
rect 5198 8186 5254 8188
rect 5278 8186 5334 8188
rect 5358 8186 5414 8188
rect 5118 8134 5164 8186
rect 5164 8134 5174 8186
rect 5198 8134 5228 8186
rect 5228 8134 5240 8186
rect 5240 8134 5254 8186
rect 5278 8134 5292 8186
rect 5292 8134 5304 8186
rect 5304 8134 5334 8186
rect 5358 8134 5368 8186
rect 5368 8134 5414 8186
rect 5118 8132 5174 8134
rect 5198 8132 5254 8134
rect 5278 8132 5334 8134
rect 5358 8132 5414 8134
rect 9833 8186 9889 8188
rect 9913 8186 9969 8188
rect 9993 8186 10049 8188
rect 10073 8186 10129 8188
rect 9833 8134 9879 8186
rect 9879 8134 9889 8186
rect 9913 8134 9943 8186
rect 9943 8134 9955 8186
rect 9955 8134 9969 8186
rect 9993 8134 10007 8186
rect 10007 8134 10019 8186
rect 10019 8134 10049 8186
rect 10073 8134 10083 8186
rect 10083 8134 10129 8186
rect 9833 8132 9889 8134
rect 9913 8132 9969 8134
rect 9993 8132 10049 8134
rect 10073 8132 10129 8134
rect 14548 8186 14604 8188
rect 14628 8186 14684 8188
rect 14708 8186 14764 8188
rect 14788 8186 14844 8188
rect 14548 8134 14594 8186
rect 14594 8134 14604 8186
rect 14628 8134 14658 8186
rect 14658 8134 14670 8186
rect 14670 8134 14684 8186
rect 14708 8134 14722 8186
rect 14722 8134 14734 8186
rect 14734 8134 14764 8186
rect 14788 8134 14798 8186
rect 14798 8134 14844 8186
rect 14548 8132 14604 8134
rect 14628 8132 14684 8134
rect 14708 8132 14764 8134
rect 14788 8132 14844 8134
rect 19263 8186 19319 8188
rect 19343 8186 19399 8188
rect 19423 8186 19479 8188
rect 19503 8186 19559 8188
rect 19263 8134 19309 8186
rect 19309 8134 19319 8186
rect 19343 8134 19373 8186
rect 19373 8134 19385 8186
rect 19385 8134 19399 8186
rect 19423 8134 19437 8186
rect 19437 8134 19449 8186
rect 19449 8134 19479 8186
rect 19503 8134 19513 8186
rect 19513 8134 19559 8186
rect 19263 8132 19319 8134
rect 19343 8132 19399 8134
rect 19423 8132 19479 8134
rect 19503 8132 19559 8134
rect 2761 7642 2817 7644
rect 2841 7642 2897 7644
rect 2921 7642 2977 7644
rect 3001 7642 3057 7644
rect 2761 7590 2807 7642
rect 2807 7590 2817 7642
rect 2841 7590 2871 7642
rect 2871 7590 2883 7642
rect 2883 7590 2897 7642
rect 2921 7590 2935 7642
rect 2935 7590 2947 7642
rect 2947 7590 2977 7642
rect 3001 7590 3011 7642
rect 3011 7590 3057 7642
rect 2761 7588 2817 7590
rect 2841 7588 2897 7590
rect 2921 7588 2977 7590
rect 3001 7588 3057 7590
rect 7476 7642 7532 7644
rect 7556 7642 7612 7644
rect 7636 7642 7692 7644
rect 7716 7642 7772 7644
rect 7476 7590 7522 7642
rect 7522 7590 7532 7642
rect 7556 7590 7586 7642
rect 7586 7590 7598 7642
rect 7598 7590 7612 7642
rect 7636 7590 7650 7642
rect 7650 7590 7662 7642
rect 7662 7590 7692 7642
rect 7716 7590 7726 7642
rect 7726 7590 7772 7642
rect 7476 7588 7532 7590
rect 7556 7588 7612 7590
rect 7636 7588 7692 7590
rect 7716 7588 7772 7590
rect 12191 7642 12247 7644
rect 12271 7642 12327 7644
rect 12351 7642 12407 7644
rect 12431 7642 12487 7644
rect 12191 7590 12237 7642
rect 12237 7590 12247 7642
rect 12271 7590 12301 7642
rect 12301 7590 12313 7642
rect 12313 7590 12327 7642
rect 12351 7590 12365 7642
rect 12365 7590 12377 7642
rect 12377 7590 12407 7642
rect 12431 7590 12441 7642
rect 12441 7590 12487 7642
rect 12191 7588 12247 7590
rect 12271 7588 12327 7590
rect 12351 7588 12407 7590
rect 12431 7588 12487 7590
rect 16906 7642 16962 7644
rect 16986 7642 17042 7644
rect 17066 7642 17122 7644
rect 17146 7642 17202 7644
rect 16906 7590 16952 7642
rect 16952 7590 16962 7642
rect 16986 7590 17016 7642
rect 17016 7590 17028 7642
rect 17028 7590 17042 7642
rect 17066 7590 17080 7642
rect 17080 7590 17092 7642
rect 17092 7590 17122 7642
rect 17146 7590 17156 7642
rect 17156 7590 17202 7642
rect 16906 7588 16962 7590
rect 16986 7588 17042 7590
rect 17066 7588 17122 7590
rect 17146 7588 17202 7590
rect 5118 7098 5174 7100
rect 5198 7098 5254 7100
rect 5278 7098 5334 7100
rect 5358 7098 5414 7100
rect 5118 7046 5164 7098
rect 5164 7046 5174 7098
rect 5198 7046 5228 7098
rect 5228 7046 5240 7098
rect 5240 7046 5254 7098
rect 5278 7046 5292 7098
rect 5292 7046 5304 7098
rect 5304 7046 5334 7098
rect 5358 7046 5368 7098
rect 5368 7046 5414 7098
rect 5118 7044 5174 7046
rect 5198 7044 5254 7046
rect 5278 7044 5334 7046
rect 5358 7044 5414 7046
rect 9833 7098 9889 7100
rect 9913 7098 9969 7100
rect 9993 7098 10049 7100
rect 10073 7098 10129 7100
rect 9833 7046 9879 7098
rect 9879 7046 9889 7098
rect 9913 7046 9943 7098
rect 9943 7046 9955 7098
rect 9955 7046 9969 7098
rect 9993 7046 10007 7098
rect 10007 7046 10019 7098
rect 10019 7046 10049 7098
rect 10073 7046 10083 7098
rect 10083 7046 10129 7098
rect 9833 7044 9889 7046
rect 9913 7044 9969 7046
rect 9993 7044 10049 7046
rect 10073 7044 10129 7046
rect 14548 7098 14604 7100
rect 14628 7098 14684 7100
rect 14708 7098 14764 7100
rect 14788 7098 14844 7100
rect 14548 7046 14594 7098
rect 14594 7046 14604 7098
rect 14628 7046 14658 7098
rect 14658 7046 14670 7098
rect 14670 7046 14684 7098
rect 14708 7046 14722 7098
rect 14722 7046 14734 7098
rect 14734 7046 14764 7098
rect 14788 7046 14798 7098
rect 14798 7046 14844 7098
rect 14548 7044 14604 7046
rect 14628 7044 14684 7046
rect 14708 7044 14764 7046
rect 14788 7044 14844 7046
rect 19263 7098 19319 7100
rect 19343 7098 19399 7100
rect 19423 7098 19479 7100
rect 19503 7098 19559 7100
rect 19263 7046 19309 7098
rect 19309 7046 19319 7098
rect 19343 7046 19373 7098
rect 19373 7046 19385 7098
rect 19385 7046 19399 7098
rect 19423 7046 19437 7098
rect 19437 7046 19449 7098
rect 19449 7046 19479 7098
rect 19503 7046 19513 7098
rect 19513 7046 19559 7098
rect 19263 7044 19319 7046
rect 19343 7044 19399 7046
rect 19423 7044 19479 7046
rect 19503 7044 19559 7046
rect 2761 6554 2817 6556
rect 2841 6554 2897 6556
rect 2921 6554 2977 6556
rect 3001 6554 3057 6556
rect 2761 6502 2807 6554
rect 2807 6502 2817 6554
rect 2841 6502 2871 6554
rect 2871 6502 2883 6554
rect 2883 6502 2897 6554
rect 2921 6502 2935 6554
rect 2935 6502 2947 6554
rect 2947 6502 2977 6554
rect 3001 6502 3011 6554
rect 3011 6502 3057 6554
rect 2761 6500 2817 6502
rect 2841 6500 2897 6502
rect 2921 6500 2977 6502
rect 3001 6500 3057 6502
rect 7476 6554 7532 6556
rect 7556 6554 7612 6556
rect 7636 6554 7692 6556
rect 7716 6554 7772 6556
rect 7476 6502 7522 6554
rect 7522 6502 7532 6554
rect 7556 6502 7586 6554
rect 7586 6502 7598 6554
rect 7598 6502 7612 6554
rect 7636 6502 7650 6554
rect 7650 6502 7662 6554
rect 7662 6502 7692 6554
rect 7716 6502 7726 6554
rect 7726 6502 7772 6554
rect 7476 6500 7532 6502
rect 7556 6500 7612 6502
rect 7636 6500 7692 6502
rect 7716 6500 7772 6502
rect 12191 6554 12247 6556
rect 12271 6554 12327 6556
rect 12351 6554 12407 6556
rect 12431 6554 12487 6556
rect 12191 6502 12237 6554
rect 12237 6502 12247 6554
rect 12271 6502 12301 6554
rect 12301 6502 12313 6554
rect 12313 6502 12327 6554
rect 12351 6502 12365 6554
rect 12365 6502 12377 6554
rect 12377 6502 12407 6554
rect 12431 6502 12441 6554
rect 12441 6502 12487 6554
rect 12191 6500 12247 6502
rect 12271 6500 12327 6502
rect 12351 6500 12407 6502
rect 12431 6500 12487 6502
rect 16906 6554 16962 6556
rect 16986 6554 17042 6556
rect 17066 6554 17122 6556
rect 17146 6554 17202 6556
rect 16906 6502 16952 6554
rect 16952 6502 16962 6554
rect 16986 6502 17016 6554
rect 17016 6502 17028 6554
rect 17028 6502 17042 6554
rect 17066 6502 17080 6554
rect 17080 6502 17092 6554
rect 17092 6502 17122 6554
rect 17146 6502 17156 6554
rect 17156 6502 17202 6554
rect 16906 6500 16962 6502
rect 16986 6500 17042 6502
rect 17066 6500 17122 6502
rect 17146 6500 17202 6502
rect 5118 6010 5174 6012
rect 5198 6010 5254 6012
rect 5278 6010 5334 6012
rect 5358 6010 5414 6012
rect 5118 5958 5164 6010
rect 5164 5958 5174 6010
rect 5198 5958 5228 6010
rect 5228 5958 5240 6010
rect 5240 5958 5254 6010
rect 5278 5958 5292 6010
rect 5292 5958 5304 6010
rect 5304 5958 5334 6010
rect 5358 5958 5368 6010
rect 5368 5958 5414 6010
rect 5118 5956 5174 5958
rect 5198 5956 5254 5958
rect 5278 5956 5334 5958
rect 5358 5956 5414 5958
rect 9833 6010 9889 6012
rect 9913 6010 9969 6012
rect 9993 6010 10049 6012
rect 10073 6010 10129 6012
rect 9833 5958 9879 6010
rect 9879 5958 9889 6010
rect 9913 5958 9943 6010
rect 9943 5958 9955 6010
rect 9955 5958 9969 6010
rect 9993 5958 10007 6010
rect 10007 5958 10019 6010
rect 10019 5958 10049 6010
rect 10073 5958 10083 6010
rect 10083 5958 10129 6010
rect 9833 5956 9889 5958
rect 9913 5956 9969 5958
rect 9993 5956 10049 5958
rect 10073 5956 10129 5958
rect 14548 6010 14604 6012
rect 14628 6010 14684 6012
rect 14708 6010 14764 6012
rect 14788 6010 14844 6012
rect 14548 5958 14594 6010
rect 14594 5958 14604 6010
rect 14628 5958 14658 6010
rect 14658 5958 14670 6010
rect 14670 5958 14684 6010
rect 14708 5958 14722 6010
rect 14722 5958 14734 6010
rect 14734 5958 14764 6010
rect 14788 5958 14798 6010
rect 14798 5958 14844 6010
rect 14548 5956 14604 5958
rect 14628 5956 14684 5958
rect 14708 5956 14764 5958
rect 14788 5956 14844 5958
rect 19263 6010 19319 6012
rect 19343 6010 19399 6012
rect 19423 6010 19479 6012
rect 19503 6010 19559 6012
rect 19263 5958 19309 6010
rect 19309 5958 19319 6010
rect 19343 5958 19373 6010
rect 19373 5958 19385 6010
rect 19385 5958 19399 6010
rect 19423 5958 19437 6010
rect 19437 5958 19449 6010
rect 19449 5958 19479 6010
rect 19503 5958 19513 6010
rect 19513 5958 19559 6010
rect 19263 5956 19319 5958
rect 19343 5956 19399 5958
rect 19423 5956 19479 5958
rect 19503 5956 19559 5958
rect 2761 5466 2817 5468
rect 2841 5466 2897 5468
rect 2921 5466 2977 5468
rect 3001 5466 3057 5468
rect 2761 5414 2807 5466
rect 2807 5414 2817 5466
rect 2841 5414 2871 5466
rect 2871 5414 2883 5466
rect 2883 5414 2897 5466
rect 2921 5414 2935 5466
rect 2935 5414 2947 5466
rect 2947 5414 2977 5466
rect 3001 5414 3011 5466
rect 3011 5414 3057 5466
rect 2761 5412 2817 5414
rect 2841 5412 2897 5414
rect 2921 5412 2977 5414
rect 3001 5412 3057 5414
rect 7476 5466 7532 5468
rect 7556 5466 7612 5468
rect 7636 5466 7692 5468
rect 7716 5466 7772 5468
rect 7476 5414 7522 5466
rect 7522 5414 7532 5466
rect 7556 5414 7586 5466
rect 7586 5414 7598 5466
rect 7598 5414 7612 5466
rect 7636 5414 7650 5466
rect 7650 5414 7662 5466
rect 7662 5414 7692 5466
rect 7716 5414 7726 5466
rect 7726 5414 7772 5466
rect 7476 5412 7532 5414
rect 7556 5412 7612 5414
rect 7636 5412 7692 5414
rect 7716 5412 7772 5414
rect 12191 5466 12247 5468
rect 12271 5466 12327 5468
rect 12351 5466 12407 5468
rect 12431 5466 12487 5468
rect 12191 5414 12237 5466
rect 12237 5414 12247 5466
rect 12271 5414 12301 5466
rect 12301 5414 12313 5466
rect 12313 5414 12327 5466
rect 12351 5414 12365 5466
rect 12365 5414 12377 5466
rect 12377 5414 12407 5466
rect 12431 5414 12441 5466
rect 12441 5414 12487 5466
rect 12191 5412 12247 5414
rect 12271 5412 12327 5414
rect 12351 5412 12407 5414
rect 12431 5412 12487 5414
rect 16906 5466 16962 5468
rect 16986 5466 17042 5468
rect 17066 5466 17122 5468
rect 17146 5466 17202 5468
rect 16906 5414 16952 5466
rect 16952 5414 16962 5466
rect 16986 5414 17016 5466
rect 17016 5414 17028 5466
rect 17028 5414 17042 5466
rect 17066 5414 17080 5466
rect 17080 5414 17092 5466
rect 17092 5414 17122 5466
rect 17146 5414 17156 5466
rect 17156 5414 17202 5466
rect 16906 5412 16962 5414
rect 16986 5412 17042 5414
rect 17066 5412 17122 5414
rect 17146 5412 17202 5414
rect 5118 4922 5174 4924
rect 5198 4922 5254 4924
rect 5278 4922 5334 4924
rect 5358 4922 5414 4924
rect 5118 4870 5164 4922
rect 5164 4870 5174 4922
rect 5198 4870 5228 4922
rect 5228 4870 5240 4922
rect 5240 4870 5254 4922
rect 5278 4870 5292 4922
rect 5292 4870 5304 4922
rect 5304 4870 5334 4922
rect 5358 4870 5368 4922
rect 5368 4870 5414 4922
rect 5118 4868 5174 4870
rect 5198 4868 5254 4870
rect 5278 4868 5334 4870
rect 5358 4868 5414 4870
rect 9833 4922 9889 4924
rect 9913 4922 9969 4924
rect 9993 4922 10049 4924
rect 10073 4922 10129 4924
rect 9833 4870 9879 4922
rect 9879 4870 9889 4922
rect 9913 4870 9943 4922
rect 9943 4870 9955 4922
rect 9955 4870 9969 4922
rect 9993 4870 10007 4922
rect 10007 4870 10019 4922
rect 10019 4870 10049 4922
rect 10073 4870 10083 4922
rect 10083 4870 10129 4922
rect 9833 4868 9889 4870
rect 9913 4868 9969 4870
rect 9993 4868 10049 4870
rect 10073 4868 10129 4870
rect 14548 4922 14604 4924
rect 14628 4922 14684 4924
rect 14708 4922 14764 4924
rect 14788 4922 14844 4924
rect 14548 4870 14594 4922
rect 14594 4870 14604 4922
rect 14628 4870 14658 4922
rect 14658 4870 14670 4922
rect 14670 4870 14684 4922
rect 14708 4870 14722 4922
rect 14722 4870 14734 4922
rect 14734 4870 14764 4922
rect 14788 4870 14798 4922
rect 14798 4870 14844 4922
rect 14548 4868 14604 4870
rect 14628 4868 14684 4870
rect 14708 4868 14764 4870
rect 14788 4868 14844 4870
rect 19263 4922 19319 4924
rect 19343 4922 19399 4924
rect 19423 4922 19479 4924
rect 19503 4922 19559 4924
rect 19263 4870 19309 4922
rect 19309 4870 19319 4922
rect 19343 4870 19373 4922
rect 19373 4870 19385 4922
rect 19385 4870 19399 4922
rect 19423 4870 19437 4922
rect 19437 4870 19449 4922
rect 19449 4870 19479 4922
rect 19503 4870 19513 4922
rect 19513 4870 19559 4922
rect 19263 4868 19319 4870
rect 19343 4868 19399 4870
rect 19423 4868 19479 4870
rect 19503 4868 19559 4870
rect 2761 4378 2817 4380
rect 2841 4378 2897 4380
rect 2921 4378 2977 4380
rect 3001 4378 3057 4380
rect 2761 4326 2807 4378
rect 2807 4326 2817 4378
rect 2841 4326 2871 4378
rect 2871 4326 2883 4378
rect 2883 4326 2897 4378
rect 2921 4326 2935 4378
rect 2935 4326 2947 4378
rect 2947 4326 2977 4378
rect 3001 4326 3011 4378
rect 3011 4326 3057 4378
rect 2761 4324 2817 4326
rect 2841 4324 2897 4326
rect 2921 4324 2977 4326
rect 3001 4324 3057 4326
rect 7476 4378 7532 4380
rect 7556 4378 7612 4380
rect 7636 4378 7692 4380
rect 7716 4378 7772 4380
rect 7476 4326 7522 4378
rect 7522 4326 7532 4378
rect 7556 4326 7586 4378
rect 7586 4326 7598 4378
rect 7598 4326 7612 4378
rect 7636 4326 7650 4378
rect 7650 4326 7662 4378
rect 7662 4326 7692 4378
rect 7716 4326 7726 4378
rect 7726 4326 7772 4378
rect 7476 4324 7532 4326
rect 7556 4324 7612 4326
rect 7636 4324 7692 4326
rect 7716 4324 7772 4326
rect 12191 4378 12247 4380
rect 12271 4378 12327 4380
rect 12351 4378 12407 4380
rect 12431 4378 12487 4380
rect 12191 4326 12237 4378
rect 12237 4326 12247 4378
rect 12271 4326 12301 4378
rect 12301 4326 12313 4378
rect 12313 4326 12327 4378
rect 12351 4326 12365 4378
rect 12365 4326 12377 4378
rect 12377 4326 12407 4378
rect 12431 4326 12441 4378
rect 12441 4326 12487 4378
rect 12191 4324 12247 4326
rect 12271 4324 12327 4326
rect 12351 4324 12407 4326
rect 12431 4324 12487 4326
rect 16906 4378 16962 4380
rect 16986 4378 17042 4380
rect 17066 4378 17122 4380
rect 17146 4378 17202 4380
rect 16906 4326 16952 4378
rect 16952 4326 16962 4378
rect 16986 4326 17016 4378
rect 17016 4326 17028 4378
rect 17028 4326 17042 4378
rect 17066 4326 17080 4378
rect 17080 4326 17092 4378
rect 17092 4326 17122 4378
rect 17146 4326 17156 4378
rect 17156 4326 17202 4378
rect 16906 4324 16962 4326
rect 16986 4324 17042 4326
rect 17066 4324 17122 4326
rect 17146 4324 17202 4326
rect 5118 3834 5174 3836
rect 5198 3834 5254 3836
rect 5278 3834 5334 3836
rect 5358 3834 5414 3836
rect 5118 3782 5164 3834
rect 5164 3782 5174 3834
rect 5198 3782 5228 3834
rect 5228 3782 5240 3834
rect 5240 3782 5254 3834
rect 5278 3782 5292 3834
rect 5292 3782 5304 3834
rect 5304 3782 5334 3834
rect 5358 3782 5368 3834
rect 5368 3782 5414 3834
rect 5118 3780 5174 3782
rect 5198 3780 5254 3782
rect 5278 3780 5334 3782
rect 5358 3780 5414 3782
rect 9833 3834 9889 3836
rect 9913 3834 9969 3836
rect 9993 3834 10049 3836
rect 10073 3834 10129 3836
rect 9833 3782 9879 3834
rect 9879 3782 9889 3834
rect 9913 3782 9943 3834
rect 9943 3782 9955 3834
rect 9955 3782 9969 3834
rect 9993 3782 10007 3834
rect 10007 3782 10019 3834
rect 10019 3782 10049 3834
rect 10073 3782 10083 3834
rect 10083 3782 10129 3834
rect 9833 3780 9889 3782
rect 9913 3780 9969 3782
rect 9993 3780 10049 3782
rect 10073 3780 10129 3782
rect 14548 3834 14604 3836
rect 14628 3834 14684 3836
rect 14708 3834 14764 3836
rect 14788 3834 14844 3836
rect 14548 3782 14594 3834
rect 14594 3782 14604 3834
rect 14628 3782 14658 3834
rect 14658 3782 14670 3834
rect 14670 3782 14684 3834
rect 14708 3782 14722 3834
rect 14722 3782 14734 3834
rect 14734 3782 14764 3834
rect 14788 3782 14798 3834
rect 14798 3782 14844 3834
rect 14548 3780 14604 3782
rect 14628 3780 14684 3782
rect 14708 3780 14764 3782
rect 14788 3780 14844 3782
rect 19263 3834 19319 3836
rect 19343 3834 19399 3836
rect 19423 3834 19479 3836
rect 19503 3834 19559 3836
rect 19263 3782 19309 3834
rect 19309 3782 19319 3834
rect 19343 3782 19373 3834
rect 19373 3782 19385 3834
rect 19385 3782 19399 3834
rect 19423 3782 19437 3834
rect 19437 3782 19449 3834
rect 19449 3782 19479 3834
rect 19503 3782 19513 3834
rect 19513 3782 19559 3834
rect 19263 3780 19319 3782
rect 19343 3780 19399 3782
rect 19423 3780 19479 3782
rect 19503 3780 19559 3782
rect 2761 3290 2817 3292
rect 2841 3290 2897 3292
rect 2921 3290 2977 3292
rect 3001 3290 3057 3292
rect 2761 3238 2807 3290
rect 2807 3238 2817 3290
rect 2841 3238 2871 3290
rect 2871 3238 2883 3290
rect 2883 3238 2897 3290
rect 2921 3238 2935 3290
rect 2935 3238 2947 3290
rect 2947 3238 2977 3290
rect 3001 3238 3011 3290
rect 3011 3238 3057 3290
rect 2761 3236 2817 3238
rect 2841 3236 2897 3238
rect 2921 3236 2977 3238
rect 3001 3236 3057 3238
rect 7476 3290 7532 3292
rect 7556 3290 7612 3292
rect 7636 3290 7692 3292
rect 7716 3290 7772 3292
rect 7476 3238 7522 3290
rect 7522 3238 7532 3290
rect 7556 3238 7586 3290
rect 7586 3238 7598 3290
rect 7598 3238 7612 3290
rect 7636 3238 7650 3290
rect 7650 3238 7662 3290
rect 7662 3238 7692 3290
rect 7716 3238 7726 3290
rect 7726 3238 7772 3290
rect 7476 3236 7532 3238
rect 7556 3236 7612 3238
rect 7636 3236 7692 3238
rect 7716 3236 7772 3238
rect 12191 3290 12247 3292
rect 12271 3290 12327 3292
rect 12351 3290 12407 3292
rect 12431 3290 12487 3292
rect 12191 3238 12237 3290
rect 12237 3238 12247 3290
rect 12271 3238 12301 3290
rect 12301 3238 12313 3290
rect 12313 3238 12327 3290
rect 12351 3238 12365 3290
rect 12365 3238 12377 3290
rect 12377 3238 12407 3290
rect 12431 3238 12441 3290
rect 12441 3238 12487 3290
rect 12191 3236 12247 3238
rect 12271 3236 12327 3238
rect 12351 3236 12407 3238
rect 12431 3236 12487 3238
rect 16906 3290 16962 3292
rect 16986 3290 17042 3292
rect 17066 3290 17122 3292
rect 17146 3290 17202 3292
rect 16906 3238 16952 3290
rect 16952 3238 16962 3290
rect 16986 3238 17016 3290
rect 17016 3238 17028 3290
rect 17028 3238 17042 3290
rect 17066 3238 17080 3290
rect 17080 3238 17092 3290
rect 17092 3238 17122 3290
rect 17146 3238 17156 3290
rect 17156 3238 17202 3290
rect 16906 3236 16962 3238
rect 16986 3236 17042 3238
rect 17066 3236 17122 3238
rect 17146 3236 17202 3238
rect 5118 2746 5174 2748
rect 5198 2746 5254 2748
rect 5278 2746 5334 2748
rect 5358 2746 5414 2748
rect 5118 2694 5164 2746
rect 5164 2694 5174 2746
rect 5198 2694 5228 2746
rect 5228 2694 5240 2746
rect 5240 2694 5254 2746
rect 5278 2694 5292 2746
rect 5292 2694 5304 2746
rect 5304 2694 5334 2746
rect 5358 2694 5368 2746
rect 5368 2694 5414 2746
rect 5118 2692 5174 2694
rect 5198 2692 5254 2694
rect 5278 2692 5334 2694
rect 5358 2692 5414 2694
rect 9833 2746 9889 2748
rect 9913 2746 9969 2748
rect 9993 2746 10049 2748
rect 10073 2746 10129 2748
rect 9833 2694 9879 2746
rect 9879 2694 9889 2746
rect 9913 2694 9943 2746
rect 9943 2694 9955 2746
rect 9955 2694 9969 2746
rect 9993 2694 10007 2746
rect 10007 2694 10019 2746
rect 10019 2694 10049 2746
rect 10073 2694 10083 2746
rect 10083 2694 10129 2746
rect 9833 2692 9889 2694
rect 9913 2692 9969 2694
rect 9993 2692 10049 2694
rect 10073 2692 10129 2694
rect 14548 2746 14604 2748
rect 14628 2746 14684 2748
rect 14708 2746 14764 2748
rect 14788 2746 14844 2748
rect 14548 2694 14594 2746
rect 14594 2694 14604 2746
rect 14628 2694 14658 2746
rect 14658 2694 14670 2746
rect 14670 2694 14684 2746
rect 14708 2694 14722 2746
rect 14722 2694 14734 2746
rect 14734 2694 14764 2746
rect 14788 2694 14798 2746
rect 14798 2694 14844 2746
rect 14548 2692 14604 2694
rect 14628 2692 14684 2694
rect 14708 2692 14764 2694
rect 14788 2692 14844 2694
rect 19263 2746 19319 2748
rect 19343 2746 19399 2748
rect 19423 2746 19479 2748
rect 19503 2746 19559 2748
rect 19263 2694 19309 2746
rect 19309 2694 19319 2746
rect 19343 2694 19373 2746
rect 19373 2694 19385 2746
rect 19385 2694 19399 2746
rect 19423 2694 19437 2746
rect 19437 2694 19449 2746
rect 19449 2694 19479 2746
rect 19503 2694 19513 2746
rect 19513 2694 19559 2746
rect 19263 2692 19319 2694
rect 19343 2692 19399 2694
rect 19423 2692 19479 2694
rect 19503 2692 19559 2694
rect 2761 2202 2817 2204
rect 2841 2202 2897 2204
rect 2921 2202 2977 2204
rect 3001 2202 3057 2204
rect 2761 2150 2807 2202
rect 2807 2150 2817 2202
rect 2841 2150 2871 2202
rect 2871 2150 2883 2202
rect 2883 2150 2897 2202
rect 2921 2150 2935 2202
rect 2935 2150 2947 2202
rect 2947 2150 2977 2202
rect 3001 2150 3011 2202
rect 3011 2150 3057 2202
rect 2761 2148 2817 2150
rect 2841 2148 2897 2150
rect 2921 2148 2977 2150
rect 3001 2148 3057 2150
rect 7476 2202 7532 2204
rect 7556 2202 7612 2204
rect 7636 2202 7692 2204
rect 7716 2202 7772 2204
rect 7476 2150 7522 2202
rect 7522 2150 7532 2202
rect 7556 2150 7586 2202
rect 7586 2150 7598 2202
rect 7598 2150 7612 2202
rect 7636 2150 7650 2202
rect 7650 2150 7662 2202
rect 7662 2150 7692 2202
rect 7716 2150 7726 2202
rect 7726 2150 7772 2202
rect 7476 2148 7532 2150
rect 7556 2148 7612 2150
rect 7636 2148 7692 2150
rect 7716 2148 7772 2150
rect 12191 2202 12247 2204
rect 12271 2202 12327 2204
rect 12351 2202 12407 2204
rect 12431 2202 12487 2204
rect 12191 2150 12237 2202
rect 12237 2150 12247 2202
rect 12271 2150 12301 2202
rect 12301 2150 12313 2202
rect 12313 2150 12327 2202
rect 12351 2150 12365 2202
rect 12365 2150 12377 2202
rect 12377 2150 12407 2202
rect 12431 2150 12441 2202
rect 12441 2150 12487 2202
rect 12191 2148 12247 2150
rect 12271 2148 12327 2150
rect 12351 2148 12407 2150
rect 12431 2148 12487 2150
rect 16906 2202 16962 2204
rect 16986 2202 17042 2204
rect 17066 2202 17122 2204
rect 17146 2202 17202 2204
rect 16906 2150 16952 2202
rect 16952 2150 16962 2202
rect 16986 2150 17016 2202
rect 17016 2150 17028 2202
rect 17028 2150 17042 2202
rect 17066 2150 17080 2202
rect 17080 2150 17092 2202
rect 17092 2150 17122 2202
rect 17146 2150 17156 2202
rect 17156 2150 17202 2202
rect 16906 2148 16962 2150
rect 16986 2148 17042 2150
rect 17066 2148 17122 2150
rect 17146 2148 17202 2150
rect 5118 1658 5174 1660
rect 5198 1658 5254 1660
rect 5278 1658 5334 1660
rect 5358 1658 5414 1660
rect 5118 1606 5164 1658
rect 5164 1606 5174 1658
rect 5198 1606 5228 1658
rect 5228 1606 5240 1658
rect 5240 1606 5254 1658
rect 5278 1606 5292 1658
rect 5292 1606 5304 1658
rect 5304 1606 5334 1658
rect 5358 1606 5368 1658
rect 5368 1606 5414 1658
rect 5118 1604 5174 1606
rect 5198 1604 5254 1606
rect 5278 1604 5334 1606
rect 5358 1604 5414 1606
rect 9833 1658 9889 1660
rect 9913 1658 9969 1660
rect 9993 1658 10049 1660
rect 10073 1658 10129 1660
rect 9833 1606 9879 1658
rect 9879 1606 9889 1658
rect 9913 1606 9943 1658
rect 9943 1606 9955 1658
rect 9955 1606 9969 1658
rect 9993 1606 10007 1658
rect 10007 1606 10019 1658
rect 10019 1606 10049 1658
rect 10073 1606 10083 1658
rect 10083 1606 10129 1658
rect 9833 1604 9889 1606
rect 9913 1604 9969 1606
rect 9993 1604 10049 1606
rect 10073 1604 10129 1606
rect 14548 1658 14604 1660
rect 14628 1658 14684 1660
rect 14708 1658 14764 1660
rect 14788 1658 14844 1660
rect 14548 1606 14594 1658
rect 14594 1606 14604 1658
rect 14628 1606 14658 1658
rect 14658 1606 14670 1658
rect 14670 1606 14684 1658
rect 14708 1606 14722 1658
rect 14722 1606 14734 1658
rect 14734 1606 14764 1658
rect 14788 1606 14798 1658
rect 14798 1606 14844 1658
rect 14548 1604 14604 1606
rect 14628 1604 14684 1606
rect 14708 1604 14764 1606
rect 14788 1604 14844 1606
rect 19263 1658 19319 1660
rect 19343 1658 19399 1660
rect 19423 1658 19479 1660
rect 19503 1658 19559 1660
rect 19263 1606 19309 1658
rect 19309 1606 19319 1658
rect 19343 1606 19373 1658
rect 19373 1606 19385 1658
rect 19385 1606 19399 1658
rect 19423 1606 19437 1658
rect 19437 1606 19449 1658
rect 19449 1606 19479 1658
rect 19503 1606 19513 1658
rect 19513 1606 19559 1658
rect 19263 1604 19319 1606
rect 19343 1604 19399 1606
rect 19423 1604 19479 1606
rect 19503 1604 19559 1606
rect 2761 1114 2817 1116
rect 2841 1114 2897 1116
rect 2921 1114 2977 1116
rect 3001 1114 3057 1116
rect 2761 1062 2807 1114
rect 2807 1062 2817 1114
rect 2841 1062 2871 1114
rect 2871 1062 2883 1114
rect 2883 1062 2897 1114
rect 2921 1062 2935 1114
rect 2935 1062 2947 1114
rect 2947 1062 2977 1114
rect 3001 1062 3011 1114
rect 3011 1062 3057 1114
rect 2761 1060 2817 1062
rect 2841 1060 2897 1062
rect 2921 1060 2977 1062
rect 3001 1060 3057 1062
rect 7476 1114 7532 1116
rect 7556 1114 7612 1116
rect 7636 1114 7692 1116
rect 7716 1114 7772 1116
rect 7476 1062 7522 1114
rect 7522 1062 7532 1114
rect 7556 1062 7586 1114
rect 7586 1062 7598 1114
rect 7598 1062 7612 1114
rect 7636 1062 7650 1114
rect 7650 1062 7662 1114
rect 7662 1062 7692 1114
rect 7716 1062 7726 1114
rect 7726 1062 7772 1114
rect 7476 1060 7532 1062
rect 7556 1060 7612 1062
rect 7636 1060 7692 1062
rect 7716 1060 7772 1062
rect 12191 1114 12247 1116
rect 12271 1114 12327 1116
rect 12351 1114 12407 1116
rect 12431 1114 12487 1116
rect 12191 1062 12237 1114
rect 12237 1062 12247 1114
rect 12271 1062 12301 1114
rect 12301 1062 12313 1114
rect 12313 1062 12327 1114
rect 12351 1062 12365 1114
rect 12365 1062 12377 1114
rect 12377 1062 12407 1114
rect 12431 1062 12441 1114
rect 12441 1062 12487 1114
rect 12191 1060 12247 1062
rect 12271 1060 12327 1062
rect 12351 1060 12407 1062
rect 12431 1060 12487 1062
rect 16906 1114 16962 1116
rect 16986 1114 17042 1116
rect 17066 1114 17122 1116
rect 17146 1114 17202 1116
rect 16906 1062 16952 1114
rect 16952 1062 16962 1114
rect 16986 1062 17016 1114
rect 17016 1062 17028 1114
rect 17028 1062 17042 1114
rect 17066 1062 17080 1114
rect 17080 1062 17092 1114
rect 17092 1062 17122 1114
rect 17146 1062 17156 1114
rect 17156 1062 17202 1114
rect 16906 1060 16962 1062
rect 16986 1060 17042 1062
rect 17066 1060 17122 1062
rect 17146 1060 17202 1062
rect 5118 570 5174 572
rect 5198 570 5254 572
rect 5278 570 5334 572
rect 5358 570 5414 572
rect 5118 518 5164 570
rect 5164 518 5174 570
rect 5198 518 5228 570
rect 5228 518 5240 570
rect 5240 518 5254 570
rect 5278 518 5292 570
rect 5292 518 5304 570
rect 5304 518 5334 570
rect 5358 518 5368 570
rect 5368 518 5414 570
rect 5118 516 5174 518
rect 5198 516 5254 518
rect 5278 516 5334 518
rect 5358 516 5414 518
rect 9833 570 9889 572
rect 9913 570 9969 572
rect 9993 570 10049 572
rect 10073 570 10129 572
rect 9833 518 9879 570
rect 9879 518 9889 570
rect 9913 518 9943 570
rect 9943 518 9955 570
rect 9955 518 9969 570
rect 9993 518 10007 570
rect 10007 518 10019 570
rect 10019 518 10049 570
rect 10073 518 10083 570
rect 10083 518 10129 570
rect 9833 516 9889 518
rect 9913 516 9969 518
rect 9993 516 10049 518
rect 10073 516 10129 518
rect 14548 570 14604 572
rect 14628 570 14684 572
rect 14708 570 14764 572
rect 14788 570 14844 572
rect 14548 518 14594 570
rect 14594 518 14604 570
rect 14628 518 14658 570
rect 14658 518 14670 570
rect 14670 518 14684 570
rect 14708 518 14722 570
rect 14722 518 14734 570
rect 14734 518 14764 570
rect 14788 518 14798 570
rect 14798 518 14844 570
rect 14548 516 14604 518
rect 14628 516 14684 518
rect 14708 516 14764 518
rect 14788 516 14844 518
rect 19263 570 19319 572
rect 19343 570 19399 572
rect 19423 570 19479 572
rect 19503 570 19559 572
rect 19263 518 19309 570
rect 19309 518 19319 570
rect 19343 518 19373 570
rect 19373 518 19385 570
rect 19385 518 19399 570
rect 19423 518 19437 570
rect 19437 518 19449 570
rect 19449 518 19479 570
rect 19503 518 19513 570
rect 19513 518 19559 570
rect 19263 516 19319 518
rect 19343 516 19399 518
rect 19423 516 19479 518
rect 19503 516 19559 518
<< metal3 >>
rect 5108 19072 5424 19073
rect 5108 19008 5114 19072
rect 5178 19008 5194 19072
rect 5258 19008 5274 19072
rect 5338 19008 5354 19072
rect 5418 19008 5424 19072
rect 5108 19007 5424 19008
rect 9823 19072 10139 19073
rect 9823 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10069 19072
rect 10133 19008 10139 19072
rect 9823 19007 10139 19008
rect 14538 19072 14854 19073
rect 14538 19008 14544 19072
rect 14608 19008 14624 19072
rect 14688 19008 14704 19072
rect 14768 19008 14784 19072
rect 14848 19008 14854 19072
rect 14538 19007 14854 19008
rect 19253 19072 19569 19073
rect 19253 19008 19259 19072
rect 19323 19008 19339 19072
rect 19403 19008 19419 19072
rect 19483 19008 19499 19072
rect 19563 19008 19569 19072
rect 19253 19007 19569 19008
rect 2751 18528 3067 18529
rect 2751 18464 2757 18528
rect 2821 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3067 18528
rect 2751 18463 3067 18464
rect 7466 18528 7782 18529
rect 7466 18464 7472 18528
rect 7536 18464 7552 18528
rect 7616 18464 7632 18528
rect 7696 18464 7712 18528
rect 7776 18464 7782 18528
rect 7466 18463 7782 18464
rect 12181 18528 12497 18529
rect 12181 18464 12187 18528
rect 12251 18464 12267 18528
rect 12331 18464 12347 18528
rect 12411 18464 12427 18528
rect 12491 18464 12497 18528
rect 12181 18463 12497 18464
rect 16896 18528 17212 18529
rect 16896 18464 16902 18528
rect 16966 18464 16982 18528
rect 17046 18464 17062 18528
rect 17126 18464 17142 18528
rect 17206 18464 17212 18528
rect 16896 18463 17212 18464
rect 5108 17984 5424 17985
rect 5108 17920 5114 17984
rect 5178 17920 5194 17984
rect 5258 17920 5274 17984
rect 5338 17920 5354 17984
rect 5418 17920 5424 17984
rect 5108 17919 5424 17920
rect 9823 17984 10139 17985
rect 9823 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10069 17984
rect 10133 17920 10139 17984
rect 9823 17919 10139 17920
rect 14538 17984 14854 17985
rect 14538 17920 14544 17984
rect 14608 17920 14624 17984
rect 14688 17920 14704 17984
rect 14768 17920 14784 17984
rect 14848 17920 14854 17984
rect 14538 17919 14854 17920
rect 19253 17984 19569 17985
rect 19253 17920 19259 17984
rect 19323 17920 19339 17984
rect 19403 17920 19419 17984
rect 19483 17920 19499 17984
rect 19563 17920 19569 17984
rect 19253 17919 19569 17920
rect 2751 17440 3067 17441
rect 2751 17376 2757 17440
rect 2821 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3067 17440
rect 2751 17375 3067 17376
rect 7466 17440 7782 17441
rect 7466 17376 7472 17440
rect 7536 17376 7552 17440
rect 7616 17376 7632 17440
rect 7696 17376 7712 17440
rect 7776 17376 7782 17440
rect 7466 17375 7782 17376
rect 12181 17440 12497 17441
rect 12181 17376 12187 17440
rect 12251 17376 12267 17440
rect 12331 17376 12347 17440
rect 12411 17376 12427 17440
rect 12491 17376 12497 17440
rect 12181 17375 12497 17376
rect 16896 17440 17212 17441
rect 16896 17376 16902 17440
rect 16966 17376 16982 17440
rect 17046 17376 17062 17440
rect 17126 17376 17142 17440
rect 17206 17376 17212 17440
rect 16896 17375 17212 17376
rect 5108 16896 5424 16897
rect 5108 16832 5114 16896
rect 5178 16832 5194 16896
rect 5258 16832 5274 16896
rect 5338 16832 5354 16896
rect 5418 16832 5424 16896
rect 5108 16831 5424 16832
rect 9823 16896 10139 16897
rect 9823 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10069 16896
rect 10133 16832 10139 16896
rect 9823 16831 10139 16832
rect 14538 16896 14854 16897
rect 14538 16832 14544 16896
rect 14608 16832 14624 16896
rect 14688 16832 14704 16896
rect 14768 16832 14784 16896
rect 14848 16832 14854 16896
rect 14538 16831 14854 16832
rect 19253 16896 19569 16897
rect 19253 16832 19259 16896
rect 19323 16832 19339 16896
rect 19403 16832 19419 16896
rect 19483 16832 19499 16896
rect 19563 16832 19569 16896
rect 19253 16831 19569 16832
rect 2751 16352 3067 16353
rect 2751 16288 2757 16352
rect 2821 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3067 16352
rect 2751 16287 3067 16288
rect 7466 16352 7782 16353
rect 7466 16288 7472 16352
rect 7536 16288 7552 16352
rect 7616 16288 7632 16352
rect 7696 16288 7712 16352
rect 7776 16288 7782 16352
rect 7466 16287 7782 16288
rect 12181 16352 12497 16353
rect 12181 16288 12187 16352
rect 12251 16288 12267 16352
rect 12331 16288 12347 16352
rect 12411 16288 12427 16352
rect 12491 16288 12497 16352
rect 12181 16287 12497 16288
rect 16896 16352 17212 16353
rect 16896 16288 16902 16352
rect 16966 16288 16982 16352
rect 17046 16288 17062 16352
rect 17126 16288 17142 16352
rect 17206 16288 17212 16352
rect 16896 16287 17212 16288
rect 5108 15808 5424 15809
rect 5108 15744 5114 15808
rect 5178 15744 5194 15808
rect 5258 15744 5274 15808
rect 5338 15744 5354 15808
rect 5418 15744 5424 15808
rect 5108 15743 5424 15744
rect 9823 15808 10139 15809
rect 9823 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10069 15808
rect 10133 15744 10139 15808
rect 9823 15743 10139 15744
rect 14538 15808 14854 15809
rect 14538 15744 14544 15808
rect 14608 15744 14624 15808
rect 14688 15744 14704 15808
rect 14768 15744 14784 15808
rect 14848 15744 14854 15808
rect 14538 15743 14854 15744
rect 19253 15808 19569 15809
rect 19253 15744 19259 15808
rect 19323 15744 19339 15808
rect 19403 15744 19419 15808
rect 19483 15744 19499 15808
rect 19563 15744 19569 15808
rect 19253 15743 19569 15744
rect 2751 15264 3067 15265
rect 2751 15200 2757 15264
rect 2821 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3067 15264
rect 2751 15199 3067 15200
rect 7466 15264 7782 15265
rect 7466 15200 7472 15264
rect 7536 15200 7552 15264
rect 7616 15200 7632 15264
rect 7696 15200 7712 15264
rect 7776 15200 7782 15264
rect 7466 15199 7782 15200
rect 12181 15264 12497 15265
rect 12181 15200 12187 15264
rect 12251 15200 12267 15264
rect 12331 15200 12347 15264
rect 12411 15200 12427 15264
rect 12491 15200 12497 15264
rect 12181 15199 12497 15200
rect 16896 15264 17212 15265
rect 16896 15200 16902 15264
rect 16966 15200 16982 15264
rect 17046 15200 17062 15264
rect 17126 15200 17142 15264
rect 17206 15200 17212 15264
rect 16896 15199 17212 15200
rect 5108 14720 5424 14721
rect 5108 14656 5114 14720
rect 5178 14656 5194 14720
rect 5258 14656 5274 14720
rect 5338 14656 5354 14720
rect 5418 14656 5424 14720
rect 5108 14655 5424 14656
rect 9823 14720 10139 14721
rect 9823 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10069 14720
rect 10133 14656 10139 14720
rect 9823 14655 10139 14656
rect 14538 14720 14854 14721
rect 14538 14656 14544 14720
rect 14608 14656 14624 14720
rect 14688 14656 14704 14720
rect 14768 14656 14784 14720
rect 14848 14656 14854 14720
rect 14538 14655 14854 14656
rect 19253 14720 19569 14721
rect 19253 14656 19259 14720
rect 19323 14656 19339 14720
rect 19403 14656 19419 14720
rect 19483 14656 19499 14720
rect 19563 14656 19569 14720
rect 19253 14655 19569 14656
rect 2751 14176 3067 14177
rect 2751 14112 2757 14176
rect 2821 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3067 14176
rect 2751 14111 3067 14112
rect 7466 14176 7782 14177
rect 7466 14112 7472 14176
rect 7536 14112 7552 14176
rect 7616 14112 7632 14176
rect 7696 14112 7712 14176
rect 7776 14112 7782 14176
rect 7466 14111 7782 14112
rect 12181 14176 12497 14177
rect 12181 14112 12187 14176
rect 12251 14112 12267 14176
rect 12331 14112 12347 14176
rect 12411 14112 12427 14176
rect 12491 14112 12497 14176
rect 12181 14111 12497 14112
rect 16896 14176 17212 14177
rect 16896 14112 16902 14176
rect 16966 14112 16982 14176
rect 17046 14112 17062 14176
rect 17126 14112 17142 14176
rect 17206 14112 17212 14176
rect 16896 14111 17212 14112
rect 5108 13632 5424 13633
rect 5108 13568 5114 13632
rect 5178 13568 5194 13632
rect 5258 13568 5274 13632
rect 5338 13568 5354 13632
rect 5418 13568 5424 13632
rect 5108 13567 5424 13568
rect 9823 13632 10139 13633
rect 9823 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10069 13632
rect 10133 13568 10139 13632
rect 9823 13567 10139 13568
rect 14538 13632 14854 13633
rect 14538 13568 14544 13632
rect 14608 13568 14624 13632
rect 14688 13568 14704 13632
rect 14768 13568 14784 13632
rect 14848 13568 14854 13632
rect 14538 13567 14854 13568
rect 19253 13632 19569 13633
rect 19253 13568 19259 13632
rect 19323 13568 19339 13632
rect 19403 13568 19419 13632
rect 19483 13568 19499 13632
rect 19563 13568 19569 13632
rect 19253 13567 19569 13568
rect 2751 13088 3067 13089
rect 2751 13024 2757 13088
rect 2821 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3067 13088
rect 2751 13023 3067 13024
rect 7466 13088 7782 13089
rect 7466 13024 7472 13088
rect 7536 13024 7552 13088
rect 7616 13024 7632 13088
rect 7696 13024 7712 13088
rect 7776 13024 7782 13088
rect 7466 13023 7782 13024
rect 12181 13088 12497 13089
rect 12181 13024 12187 13088
rect 12251 13024 12267 13088
rect 12331 13024 12347 13088
rect 12411 13024 12427 13088
rect 12491 13024 12497 13088
rect 12181 13023 12497 13024
rect 16896 13088 17212 13089
rect 16896 13024 16902 13088
rect 16966 13024 16982 13088
rect 17046 13024 17062 13088
rect 17126 13024 17142 13088
rect 17206 13024 17212 13088
rect 16896 13023 17212 13024
rect 5108 12544 5424 12545
rect 5108 12480 5114 12544
rect 5178 12480 5194 12544
rect 5258 12480 5274 12544
rect 5338 12480 5354 12544
rect 5418 12480 5424 12544
rect 5108 12479 5424 12480
rect 9823 12544 10139 12545
rect 9823 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10069 12544
rect 10133 12480 10139 12544
rect 9823 12479 10139 12480
rect 14538 12544 14854 12545
rect 14538 12480 14544 12544
rect 14608 12480 14624 12544
rect 14688 12480 14704 12544
rect 14768 12480 14784 12544
rect 14848 12480 14854 12544
rect 14538 12479 14854 12480
rect 19253 12544 19569 12545
rect 19253 12480 19259 12544
rect 19323 12480 19339 12544
rect 19403 12480 19419 12544
rect 19483 12480 19499 12544
rect 19563 12480 19569 12544
rect 19253 12479 19569 12480
rect 2751 12000 3067 12001
rect 2751 11936 2757 12000
rect 2821 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3067 12000
rect 2751 11935 3067 11936
rect 7466 12000 7782 12001
rect 7466 11936 7472 12000
rect 7536 11936 7552 12000
rect 7616 11936 7632 12000
rect 7696 11936 7712 12000
rect 7776 11936 7782 12000
rect 7466 11935 7782 11936
rect 12181 12000 12497 12001
rect 12181 11936 12187 12000
rect 12251 11936 12267 12000
rect 12331 11936 12347 12000
rect 12411 11936 12427 12000
rect 12491 11936 12497 12000
rect 12181 11935 12497 11936
rect 16896 12000 17212 12001
rect 16896 11936 16902 12000
rect 16966 11936 16982 12000
rect 17046 11936 17062 12000
rect 17126 11936 17142 12000
rect 17206 11936 17212 12000
rect 16896 11935 17212 11936
rect 5108 11456 5424 11457
rect 5108 11392 5114 11456
rect 5178 11392 5194 11456
rect 5258 11392 5274 11456
rect 5338 11392 5354 11456
rect 5418 11392 5424 11456
rect 5108 11391 5424 11392
rect 9823 11456 10139 11457
rect 9823 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10069 11456
rect 10133 11392 10139 11456
rect 9823 11391 10139 11392
rect 14538 11456 14854 11457
rect 14538 11392 14544 11456
rect 14608 11392 14624 11456
rect 14688 11392 14704 11456
rect 14768 11392 14784 11456
rect 14848 11392 14854 11456
rect 14538 11391 14854 11392
rect 19253 11456 19569 11457
rect 19253 11392 19259 11456
rect 19323 11392 19339 11456
rect 19403 11392 19419 11456
rect 19483 11392 19499 11456
rect 19563 11392 19569 11456
rect 19253 11391 19569 11392
rect 2751 10912 3067 10913
rect 2751 10848 2757 10912
rect 2821 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3067 10912
rect 2751 10847 3067 10848
rect 7466 10912 7782 10913
rect 7466 10848 7472 10912
rect 7536 10848 7552 10912
rect 7616 10848 7632 10912
rect 7696 10848 7712 10912
rect 7776 10848 7782 10912
rect 7466 10847 7782 10848
rect 12181 10912 12497 10913
rect 12181 10848 12187 10912
rect 12251 10848 12267 10912
rect 12331 10848 12347 10912
rect 12411 10848 12427 10912
rect 12491 10848 12497 10912
rect 12181 10847 12497 10848
rect 16896 10912 17212 10913
rect 16896 10848 16902 10912
rect 16966 10848 16982 10912
rect 17046 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17212 10912
rect 16896 10847 17212 10848
rect 5108 10368 5424 10369
rect 5108 10304 5114 10368
rect 5178 10304 5194 10368
rect 5258 10304 5274 10368
rect 5338 10304 5354 10368
rect 5418 10304 5424 10368
rect 5108 10303 5424 10304
rect 9823 10368 10139 10369
rect 9823 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10069 10368
rect 10133 10304 10139 10368
rect 9823 10303 10139 10304
rect 14538 10368 14854 10369
rect 14538 10304 14544 10368
rect 14608 10304 14624 10368
rect 14688 10304 14704 10368
rect 14768 10304 14784 10368
rect 14848 10304 14854 10368
rect 14538 10303 14854 10304
rect 19253 10368 19569 10369
rect 19253 10304 19259 10368
rect 19323 10304 19339 10368
rect 19403 10304 19419 10368
rect 19483 10304 19499 10368
rect 19563 10304 19569 10368
rect 19253 10303 19569 10304
rect 19057 9890 19123 9893
rect 19600 9890 20000 9920
rect 19057 9888 20000 9890
rect 19057 9832 19062 9888
rect 19118 9832 20000 9888
rect 19057 9830 20000 9832
rect 19057 9827 19123 9830
rect 2751 9824 3067 9825
rect 2751 9760 2757 9824
rect 2821 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3067 9824
rect 2751 9759 3067 9760
rect 7466 9824 7782 9825
rect 7466 9760 7472 9824
rect 7536 9760 7552 9824
rect 7616 9760 7632 9824
rect 7696 9760 7712 9824
rect 7776 9760 7782 9824
rect 7466 9759 7782 9760
rect 12181 9824 12497 9825
rect 12181 9760 12187 9824
rect 12251 9760 12267 9824
rect 12331 9760 12347 9824
rect 12411 9760 12427 9824
rect 12491 9760 12497 9824
rect 12181 9759 12497 9760
rect 16896 9824 17212 9825
rect 16896 9760 16902 9824
rect 16966 9760 16982 9824
rect 17046 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17212 9824
rect 19600 9800 20000 9830
rect 16896 9759 17212 9760
rect 5108 9280 5424 9281
rect 5108 9216 5114 9280
rect 5178 9216 5194 9280
rect 5258 9216 5274 9280
rect 5338 9216 5354 9280
rect 5418 9216 5424 9280
rect 5108 9215 5424 9216
rect 9823 9280 10139 9281
rect 9823 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10069 9280
rect 10133 9216 10139 9280
rect 9823 9215 10139 9216
rect 14538 9280 14854 9281
rect 14538 9216 14544 9280
rect 14608 9216 14624 9280
rect 14688 9216 14704 9280
rect 14768 9216 14784 9280
rect 14848 9216 14854 9280
rect 14538 9215 14854 9216
rect 19253 9280 19569 9281
rect 19253 9216 19259 9280
rect 19323 9216 19339 9280
rect 19403 9216 19419 9280
rect 19483 9216 19499 9280
rect 19563 9216 19569 9280
rect 19253 9215 19569 9216
rect 2751 8736 3067 8737
rect 2751 8672 2757 8736
rect 2821 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3067 8736
rect 2751 8671 3067 8672
rect 7466 8736 7782 8737
rect 7466 8672 7472 8736
rect 7536 8672 7552 8736
rect 7616 8672 7632 8736
rect 7696 8672 7712 8736
rect 7776 8672 7782 8736
rect 7466 8671 7782 8672
rect 12181 8736 12497 8737
rect 12181 8672 12187 8736
rect 12251 8672 12267 8736
rect 12331 8672 12347 8736
rect 12411 8672 12427 8736
rect 12491 8672 12497 8736
rect 12181 8671 12497 8672
rect 16896 8736 17212 8737
rect 16896 8672 16902 8736
rect 16966 8672 16982 8736
rect 17046 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17212 8736
rect 16896 8671 17212 8672
rect 5108 8192 5424 8193
rect 5108 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5354 8192
rect 5418 8128 5424 8192
rect 5108 8127 5424 8128
rect 9823 8192 10139 8193
rect 9823 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10069 8192
rect 10133 8128 10139 8192
rect 9823 8127 10139 8128
rect 14538 8192 14854 8193
rect 14538 8128 14544 8192
rect 14608 8128 14624 8192
rect 14688 8128 14704 8192
rect 14768 8128 14784 8192
rect 14848 8128 14854 8192
rect 14538 8127 14854 8128
rect 19253 8192 19569 8193
rect 19253 8128 19259 8192
rect 19323 8128 19339 8192
rect 19403 8128 19419 8192
rect 19483 8128 19499 8192
rect 19563 8128 19569 8192
rect 19253 8127 19569 8128
rect 2751 7648 3067 7649
rect 2751 7584 2757 7648
rect 2821 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3067 7648
rect 2751 7583 3067 7584
rect 7466 7648 7782 7649
rect 7466 7584 7472 7648
rect 7536 7584 7552 7648
rect 7616 7584 7632 7648
rect 7696 7584 7712 7648
rect 7776 7584 7782 7648
rect 7466 7583 7782 7584
rect 12181 7648 12497 7649
rect 12181 7584 12187 7648
rect 12251 7584 12267 7648
rect 12331 7584 12347 7648
rect 12411 7584 12427 7648
rect 12491 7584 12497 7648
rect 12181 7583 12497 7584
rect 16896 7648 17212 7649
rect 16896 7584 16902 7648
rect 16966 7584 16982 7648
rect 17046 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17212 7648
rect 16896 7583 17212 7584
rect 5108 7104 5424 7105
rect 5108 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5354 7104
rect 5418 7040 5424 7104
rect 5108 7039 5424 7040
rect 9823 7104 10139 7105
rect 9823 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10069 7104
rect 10133 7040 10139 7104
rect 9823 7039 10139 7040
rect 14538 7104 14854 7105
rect 14538 7040 14544 7104
rect 14608 7040 14624 7104
rect 14688 7040 14704 7104
rect 14768 7040 14784 7104
rect 14848 7040 14854 7104
rect 14538 7039 14854 7040
rect 19253 7104 19569 7105
rect 19253 7040 19259 7104
rect 19323 7040 19339 7104
rect 19403 7040 19419 7104
rect 19483 7040 19499 7104
rect 19563 7040 19569 7104
rect 19253 7039 19569 7040
rect 2751 6560 3067 6561
rect 2751 6496 2757 6560
rect 2821 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3067 6560
rect 2751 6495 3067 6496
rect 7466 6560 7782 6561
rect 7466 6496 7472 6560
rect 7536 6496 7552 6560
rect 7616 6496 7632 6560
rect 7696 6496 7712 6560
rect 7776 6496 7782 6560
rect 7466 6495 7782 6496
rect 12181 6560 12497 6561
rect 12181 6496 12187 6560
rect 12251 6496 12267 6560
rect 12331 6496 12347 6560
rect 12411 6496 12427 6560
rect 12491 6496 12497 6560
rect 12181 6495 12497 6496
rect 16896 6560 17212 6561
rect 16896 6496 16902 6560
rect 16966 6496 16982 6560
rect 17046 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17212 6560
rect 16896 6495 17212 6496
rect 5108 6016 5424 6017
rect 5108 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5354 6016
rect 5418 5952 5424 6016
rect 5108 5951 5424 5952
rect 9823 6016 10139 6017
rect 9823 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10069 6016
rect 10133 5952 10139 6016
rect 9823 5951 10139 5952
rect 14538 6016 14854 6017
rect 14538 5952 14544 6016
rect 14608 5952 14624 6016
rect 14688 5952 14704 6016
rect 14768 5952 14784 6016
rect 14848 5952 14854 6016
rect 14538 5951 14854 5952
rect 19253 6016 19569 6017
rect 19253 5952 19259 6016
rect 19323 5952 19339 6016
rect 19403 5952 19419 6016
rect 19483 5952 19499 6016
rect 19563 5952 19569 6016
rect 19253 5951 19569 5952
rect 2751 5472 3067 5473
rect 2751 5408 2757 5472
rect 2821 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3067 5472
rect 2751 5407 3067 5408
rect 7466 5472 7782 5473
rect 7466 5408 7472 5472
rect 7536 5408 7552 5472
rect 7616 5408 7632 5472
rect 7696 5408 7712 5472
rect 7776 5408 7782 5472
rect 7466 5407 7782 5408
rect 12181 5472 12497 5473
rect 12181 5408 12187 5472
rect 12251 5408 12267 5472
rect 12331 5408 12347 5472
rect 12411 5408 12427 5472
rect 12491 5408 12497 5472
rect 12181 5407 12497 5408
rect 16896 5472 17212 5473
rect 16896 5408 16902 5472
rect 16966 5408 16982 5472
rect 17046 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17212 5472
rect 16896 5407 17212 5408
rect 5108 4928 5424 4929
rect 5108 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5354 4928
rect 5418 4864 5424 4928
rect 5108 4863 5424 4864
rect 9823 4928 10139 4929
rect 9823 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10069 4928
rect 10133 4864 10139 4928
rect 9823 4863 10139 4864
rect 14538 4928 14854 4929
rect 14538 4864 14544 4928
rect 14608 4864 14624 4928
rect 14688 4864 14704 4928
rect 14768 4864 14784 4928
rect 14848 4864 14854 4928
rect 14538 4863 14854 4864
rect 19253 4928 19569 4929
rect 19253 4864 19259 4928
rect 19323 4864 19339 4928
rect 19403 4864 19419 4928
rect 19483 4864 19499 4928
rect 19563 4864 19569 4928
rect 19253 4863 19569 4864
rect 2751 4384 3067 4385
rect 2751 4320 2757 4384
rect 2821 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3067 4384
rect 2751 4319 3067 4320
rect 7466 4384 7782 4385
rect 7466 4320 7472 4384
rect 7536 4320 7552 4384
rect 7616 4320 7632 4384
rect 7696 4320 7712 4384
rect 7776 4320 7782 4384
rect 7466 4319 7782 4320
rect 12181 4384 12497 4385
rect 12181 4320 12187 4384
rect 12251 4320 12267 4384
rect 12331 4320 12347 4384
rect 12411 4320 12427 4384
rect 12491 4320 12497 4384
rect 12181 4319 12497 4320
rect 16896 4384 17212 4385
rect 16896 4320 16902 4384
rect 16966 4320 16982 4384
rect 17046 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17212 4384
rect 16896 4319 17212 4320
rect 5108 3840 5424 3841
rect 5108 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5354 3840
rect 5418 3776 5424 3840
rect 5108 3775 5424 3776
rect 9823 3840 10139 3841
rect 9823 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10069 3840
rect 10133 3776 10139 3840
rect 9823 3775 10139 3776
rect 14538 3840 14854 3841
rect 14538 3776 14544 3840
rect 14608 3776 14624 3840
rect 14688 3776 14704 3840
rect 14768 3776 14784 3840
rect 14848 3776 14854 3840
rect 14538 3775 14854 3776
rect 19253 3840 19569 3841
rect 19253 3776 19259 3840
rect 19323 3776 19339 3840
rect 19403 3776 19419 3840
rect 19483 3776 19499 3840
rect 19563 3776 19569 3840
rect 19253 3775 19569 3776
rect 2751 3296 3067 3297
rect 2751 3232 2757 3296
rect 2821 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3067 3296
rect 2751 3231 3067 3232
rect 7466 3296 7782 3297
rect 7466 3232 7472 3296
rect 7536 3232 7552 3296
rect 7616 3232 7632 3296
rect 7696 3232 7712 3296
rect 7776 3232 7782 3296
rect 7466 3231 7782 3232
rect 12181 3296 12497 3297
rect 12181 3232 12187 3296
rect 12251 3232 12267 3296
rect 12331 3232 12347 3296
rect 12411 3232 12427 3296
rect 12491 3232 12497 3296
rect 12181 3231 12497 3232
rect 16896 3296 17212 3297
rect 16896 3232 16902 3296
rect 16966 3232 16982 3296
rect 17046 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17212 3296
rect 16896 3231 17212 3232
rect 5108 2752 5424 2753
rect 5108 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5354 2752
rect 5418 2688 5424 2752
rect 5108 2687 5424 2688
rect 9823 2752 10139 2753
rect 9823 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10069 2752
rect 10133 2688 10139 2752
rect 9823 2687 10139 2688
rect 14538 2752 14854 2753
rect 14538 2688 14544 2752
rect 14608 2688 14624 2752
rect 14688 2688 14704 2752
rect 14768 2688 14784 2752
rect 14848 2688 14854 2752
rect 14538 2687 14854 2688
rect 19253 2752 19569 2753
rect 19253 2688 19259 2752
rect 19323 2688 19339 2752
rect 19403 2688 19419 2752
rect 19483 2688 19499 2752
rect 19563 2688 19569 2752
rect 19253 2687 19569 2688
rect 2751 2208 3067 2209
rect 2751 2144 2757 2208
rect 2821 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3067 2208
rect 2751 2143 3067 2144
rect 7466 2208 7782 2209
rect 7466 2144 7472 2208
rect 7536 2144 7552 2208
rect 7616 2144 7632 2208
rect 7696 2144 7712 2208
rect 7776 2144 7782 2208
rect 7466 2143 7782 2144
rect 12181 2208 12497 2209
rect 12181 2144 12187 2208
rect 12251 2144 12267 2208
rect 12331 2144 12347 2208
rect 12411 2144 12427 2208
rect 12491 2144 12497 2208
rect 12181 2143 12497 2144
rect 16896 2208 17212 2209
rect 16896 2144 16902 2208
rect 16966 2144 16982 2208
rect 17046 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17212 2208
rect 16896 2143 17212 2144
rect 5108 1664 5424 1665
rect 5108 1600 5114 1664
rect 5178 1600 5194 1664
rect 5258 1600 5274 1664
rect 5338 1600 5354 1664
rect 5418 1600 5424 1664
rect 5108 1599 5424 1600
rect 9823 1664 10139 1665
rect 9823 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10069 1664
rect 10133 1600 10139 1664
rect 9823 1599 10139 1600
rect 14538 1664 14854 1665
rect 14538 1600 14544 1664
rect 14608 1600 14624 1664
rect 14688 1600 14704 1664
rect 14768 1600 14784 1664
rect 14848 1600 14854 1664
rect 14538 1599 14854 1600
rect 19253 1664 19569 1665
rect 19253 1600 19259 1664
rect 19323 1600 19339 1664
rect 19403 1600 19419 1664
rect 19483 1600 19499 1664
rect 19563 1600 19569 1664
rect 19253 1599 19569 1600
rect 2751 1120 3067 1121
rect 2751 1056 2757 1120
rect 2821 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3067 1120
rect 2751 1055 3067 1056
rect 7466 1120 7782 1121
rect 7466 1056 7472 1120
rect 7536 1056 7552 1120
rect 7616 1056 7632 1120
rect 7696 1056 7712 1120
rect 7776 1056 7782 1120
rect 7466 1055 7782 1056
rect 12181 1120 12497 1121
rect 12181 1056 12187 1120
rect 12251 1056 12267 1120
rect 12331 1056 12347 1120
rect 12411 1056 12427 1120
rect 12491 1056 12497 1120
rect 12181 1055 12497 1056
rect 16896 1120 17212 1121
rect 16896 1056 16902 1120
rect 16966 1056 16982 1120
rect 17046 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17212 1120
rect 16896 1055 17212 1056
rect 5108 576 5424 577
rect 5108 512 5114 576
rect 5178 512 5194 576
rect 5258 512 5274 576
rect 5338 512 5354 576
rect 5418 512 5424 576
rect 5108 511 5424 512
rect 9823 576 10139 577
rect 9823 512 9829 576
rect 9893 512 9909 576
rect 9973 512 9989 576
rect 10053 512 10069 576
rect 10133 512 10139 576
rect 9823 511 10139 512
rect 14538 576 14854 577
rect 14538 512 14544 576
rect 14608 512 14624 576
rect 14688 512 14704 576
rect 14768 512 14784 576
rect 14848 512 14854 576
rect 14538 511 14854 512
rect 19253 576 19569 577
rect 19253 512 19259 576
rect 19323 512 19339 576
rect 19403 512 19419 576
rect 19483 512 19499 576
rect 19563 512 19569 576
rect 19253 511 19569 512
<< via3 >>
rect 5114 19068 5178 19072
rect 5114 19012 5118 19068
rect 5118 19012 5174 19068
rect 5174 19012 5178 19068
rect 5114 19008 5178 19012
rect 5194 19068 5258 19072
rect 5194 19012 5198 19068
rect 5198 19012 5254 19068
rect 5254 19012 5258 19068
rect 5194 19008 5258 19012
rect 5274 19068 5338 19072
rect 5274 19012 5278 19068
rect 5278 19012 5334 19068
rect 5334 19012 5338 19068
rect 5274 19008 5338 19012
rect 5354 19068 5418 19072
rect 5354 19012 5358 19068
rect 5358 19012 5414 19068
rect 5414 19012 5418 19068
rect 5354 19008 5418 19012
rect 9829 19068 9893 19072
rect 9829 19012 9833 19068
rect 9833 19012 9889 19068
rect 9889 19012 9893 19068
rect 9829 19008 9893 19012
rect 9909 19068 9973 19072
rect 9909 19012 9913 19068
rect 9913 19012 9969 19068
rect 9969 19012 9973 19068
rect 9909 19008 9973 19012
rect 9989 19068 10053 19072
rect 9989 19012 9993 19068
rect 9993 19012 10049 19068
rect 10049 19012 10053 19068
rect 9989 19008 10053 19012
rect 10069 19068 10133 19072
rect 10069 19012 10073 19068
rect 10073 19012 10129 19068
rect 10129 19012 10133 19068
rect 10069 19008 10133 19012
rect 14544 19068 14608 19072
rect 14544 19012 14548 19068
rect 14548 19012 14604 19068
rect 14604 19012 14608 19068
rect 14544 19008 14608 19012
rect 14624 19068 14688 19072
rect 14624 19012 14628 19068
rect 14628 19012 14684 19068
rect 14684 19012 14688 19068
rect 14624 19008 14688 19012
rect 14704 19068 14768 19072
rect 14704 19012 14708 19068
rect 14708 19012 14764 19068
rect 14764 19012 14768 19068
rect 14704 19008 14768 19012
rect 14784 19068 14848 19072
rect 14784 19012 14788 19068
rect 14788 19012 14844 19068
rect 14844 19012 14848 19068
rect 14784 19008 14848 19012
rect 19259 19068 19323 19072
rect 19259 19012 19263 19068
rect 19263 19012 19319 19068
rect 19319 19012 19323 19068
rect 19259 19008 19323 19012
rect 19339 19068 19403 19072
rect 19339 19012 19343 19068
rect 19343 19012 19399 19068
rect 19399 19012 19403 19068
rect 19339 19008 19403 19012
rect 19419 19068 19483 19072
rect 19419 19012 19423 19068
rect 19423 19012 19479 19068
rect 19479 19012 19483 19068
rect 19419 19008 19483 19012
rect 19499 19068 19563 19072
rect 19499 19012 19503 19068
rect 19503 19012 19559 19068
rect 19559 19012 19563 19068
rect 19499 19008 19563 19012
rect 2757 18524 2821 18528
rect 2757 18468 2761 18524
rect 2761 18468 2817 18524
rect 2817 18468 2821 18524
rect 2757 18464 2821 18468
rect 2837 18524 2901 18528
rect 2837 18468 2841 18524
rect 2841 18468 2897 18524
rect 2897 18468 2901 18524
rect 2837 18464 2901 18468
rect 2917 18524 2981 18528
rect 2917 18468 2921 18524
rect 2921 18468 2977 18524
rect 2977 18468 2981 18524
rect 2917 18464 2981 18468
rect 2997 18524 3061 18528
rect 2997 18468 3001 18524
rect 3001 18468 3057 18524
rect 3057 18468 3061 18524
rect 2997 18464 3061 18468
rect 7472 18524 7536 18528
rect 7472 18468 7476 18524
rect 7476 18468 7532 18524
rect 7532 18468 7536 18524
rect 7472 18464 7536 18468
rect 7552 18524 7616 18528
rect 7552 18468 7556 18524
rect 7556 18468 7612 18524
rect 7612 18468 7616 18524
rect 7552 18464 7616 18468
rect 7632 18524 7696 18528
rect 7632 18468 7636 18524
rect 7636 18468 7692 18524
rect 7692 18468 7696 18524
rect 7632 18464 7696 18468
rect 7712 18524 7776 18528
rect 7712 18468 7716 18524
rect 7716 18468 7772 18524
rect 7772 18468 7776 18524
rect 7712 18464 7776 18468
rect 12187 18524 12251 18528
rect 12187 18468 12191 18524
rect 12191 18468 12247 18524
rect 12247 18468 12251 18524
rect 12187 18464 12251 18468
rect 12267 18524 12331 18528
rect 12267 18468 12271 18524
rect 12271 18468 12327 18524
rect 12327 18468 12331 18524
rect 12267 18464 12331 18468
rect 12347 18524 12411 18528
rect 12347 18468 12351 18524
rect 12351 18468 12407 18524
rect 12407 18468 12411 18524
rect 12347 18464 12411 18468
rect 12427 18524 12491 18528
rect 12427 18468 12431 18524
rect 12431 18468 12487 18524
rect 12487 18468 12491 18524
rect 12427 18464 12491 18468
rect 16902 18524 16966 18528
rect 16902 18468 16906 18524
rect 16906 18468 16962 18524
rect 16962 18468 16966 18524
rect 16902 18464 16966 18468
rect 16982 18524 17046 18528
rect 16982 18468 16986 18524
rect 16986 18468 17042 18524
rect 17042 18468 17046 18524
rect 16982 18464 17046 18468
rect 17062 18524 17126 18528
rect 17062 18468 17066 18524
rect 17066 18468 17122 18524
rect 17122 18468 17126 18524
rect 17062 18464 17126 18468
rect 17142 18524 17206 18528
rect 17142 18468 17146 18524
rect 17146 18468 17202 18524
rect 17202 18468 17206 18524
rect 17142 18464 17206 18468
rect 5114 17980 5178 17984
rect 5114 17924 5118 17980
rect 5118 17924 5174 17980
rect 5174 17924 5178 17980
rect 5114 17920 5178 17924
rect 5194 17980 5258 17984
rect 5194 17924 5198 17980
rect 5198 17924 5254 17980
rect 5254 17924 5258 17980
rect 5194 17920 5258 17924
rect 5274 17980 5338 17984
rect 5274 17924 5278 17980
rect 5278 17924 5334 17980
rect 5334 17924 5338 17980
rect 5274 17920 5338 17924
rect 5354 17980 5418 17984
rect 5354 17924 5358 17980
rect 5358 17924 5414 17980
rect 5414 17924 5418 17980
rect 5354 17920 5418 17924
rect 9829 17980 9893 17984
rect 9829 17924 9833 17980
rect 9833 17924 9889 17980
rect 9889 17924 9893 17980
rect 9829 17920 9893 17924
rect 9909 17980 9973 17984
rect 9909 17924 9913 17980
rect 9913 17924 9969 17980
rect 9969 17924 9973 17980
rect 9909 17920 9973 17924
rect 9989 17980 10053 17984
rect 9989 17924 9993 17980
rect 9993 17924 10049 17980
rect 10049 17924 10053 17980
rect 9989 17920 10053 17924
rect 10069 17980 10133 17984
rect 10069 17924 10073 17980
rect 10073 17924 10129 17980
rect 10129 17924 10133 17980
rect 10069 17920 10133 17924
rect 14544 17980 14608 17984
rect 14544 17924 14548 17980
rect 14548 17924 14604 17980
rect 14604 17924 14608 17980
rect 14544 17920 14608 17924
rect 14624 17980 14688 17984
rect 14624 17924 14628 17980
rect 14628 17924 14684 17980
rect 14684 17924 14688 17980
rect 14624 17920 14688 17924
rect 14704 17980 14768 17984
rect 14704 17924 14708 17980
rect 14708 17924 14764 17980
rect 14764 17924 14768 17980
rect 14704 17920 14768 17924
rect 14784 17980 14848 17984
rect 14784 17924 14788 17980
rect 14788 17924 14844 17980
rect 14844 17924 14848 17980
rect 14784 17920 14848 17924
rect 19259 17980 19323 17984
rect 19259 17924 19263 17980
rect 19263 17924 19319 17980
rect 19319 17924 19323 17980
rect 19259 17920 19323 17924
rect 19339 17980 19403 17984
rect 19339 17924 19343 17980
rect 19343 17924 19399 17980
rect 19399 17924 19403 17980
rect 19339 17920 19403 17924
rect 19419 17980 19483 17984
rect 19419 17924 19423 17980
rect 19423 17924 19479 17980
rect 19479 17924 19483 17980
rect 19419 17920 19483 17924
rect 19499 17980 19563 17984
rect 19499 17924 19503 17980
rect 19503 17924 19559 17980
rect 19559 17924 19563 17980
rect 19499 17920 19563 17924
rect 2757 17436 2821 17440
rect 2757 17380 2761 17436
rect 2761 17380 2817 17436
rect 2817 17380 2821 17436
rect 2757 17376 2821 17380
rect 2837 17436 2901 17440
rect 2837 17380 2841 17436
rect 2841 17380 2897 17436
rect 2897 17380 2901 17436
rect 2837 17376 2901 17380
rect 2917 17436 2981 17440
rect 2917 17380 2921 17436
rect 2921 17380 2977 17436
rect 2977 17380 2981 17436
rect 2917 17376 2981 17380
rect 2997 17436 3061 17440
rect 2997 17380 3001 17436
rect 3001 17380 3057 17436
rect 3057 17380 3061 17436
rect 2997 17376 3061 17380
rect 7472 17436 7536 17440
rect 7472 17380 7476 17436
rect 7476 17380 7532 17436
rect 7532 17380 7536 17436
rect 7472 17376 7536 17380
rect 7552 17436 7616 17440
rect 7552 17380 7556 17436
rect 7556 17380 7612 17436
rect 7612 17380 7616 17436
rect 7552 17376 7616 17380
rect 7632 17436 7696 17440
rect 7632 17380 7636 17436
rect 7636 17380 7692 17436
rect 7692 17380 7696 17436
rect 7632 17376 7696 17380
rect 7712 17436 7776 17440
rect 7712 17380 7716 17436
rect 7716 17380 7772 17436
rect 7772 17380 7776 17436
rect 7712 17376 7776 17380
rect 12187 17436 12251 17440
rect 12187 17380 12191 17436
rect 12191 17380 12247 17436
rect 12247 17380 12251 17436
rect 12187 17376 12251 17380
rect 12267 17436 12331 17440
rect 12267 17380 12271 17436
rect 12271 17380 12327 17436
rect 12327 17380 12331 17436
rect 12267 17376 12331 17380
rect 12347 17436 12411 17440
rect 12347 17380 12351 17436
rect 12351 17380 12407 17436
rect 12407 17380 12411 17436
rect 12347 17376 12411 17380
rect 12427 17436 12491 17440
rect 12427 17380 12431 17436
rect 12431 17380 12487 17436
rect 12487 17380 12491 17436
rect 12427 17376 12491 17380
rect 16902 17436 16966 17440
rect 16902 17380 16906 17436
rect 16906 17380 16962 17436
rect 16962 17380 16966 17436
rect 16902 17376 16966 17380
rect 16982 17436 17046 17440
rect 16982 17380 16986 17436
rect 16986 17380 17042 17436
rect 17042 17380 17046 17436
rect 16982 17376 17046 17380
rect 17062 17436 17126 17440
rect 17062 17380 17066 17436
rect 17066 17380 17122 17436
rect 17122 17380 17126 17436
rect 17062 17376 17126 17380
rect 17142 17436 17206 17440
rect 17142 17380 17146 17436
rect 17146 17380 17202 17436
rect 17202 17380 17206 17436
rect 17142 17376 17206 17380
rect 5114 16892 5178 16896
rect 5114 16836 5118 16892
rect 5118 16836 5174 16892
rect 5174 16836 5178 16892
rect 5114 16832 5178 16836
rect 5194 16892 5258 16896
rect 5194 16836 5198 16892
rect 5198 16836 5254 16892
rect 5254 16836 5258 16892
rect 5194 16832 5258 16836
rect 5274 16892 5338 16896
rect 5274 16836 5278 16892
rect 5278 16836 5334 16892
rect 5334 16836 5338 16892
rect 5274 16832 5338 16836
rect 5354 16892 5418 16896
rect 5354 16836 5358 16892
rect 5358 16836 5414 16892
rect 5414 16836 5418 16892
rect 5354 16832 5418 16836
rect 9829 16892 9893 16896
rect 9829 16836 9833 16892
rect 9833 16836 9889 16892
rect 9889 16836 9893 16892
rect 9829 16832 9893 16836
rect 9909 16892 9973 16896
rect 9909 16836 9913 16892
rect 9913 16836 9969 16892
rect 9969 16836 9973 16892
rect 9909 16832 9973 16836
rect 9989 16892 10053 16896
rect 9989 16836 9993 16892
rect 9993 16836 10049 16892
rect 10049 16836 10053 16892
rect 9989 16832 10053 16836
rect 10069 16892 10133 16896
rect 10069 16836 10073 16892
rect 10073 16836 10129 16892
rect 10129 16836 10133 16892
rect 10069 16832 10133 16836
rect 14544 16892 14608 16896
rect 14544 16836 14548 16892
rect 14548 16836 14604 16892
rect 14604 16836 14608 16892
rect 14544 16832 14608 16836
rect 14624 16892 14688 16896
rect 14624 16836 14628 16892
rect 14628 16836 14684 16892
rect 14684 16836 14688 16892
rect 14624 16832 14688 16836
rect 14704 16892 14768 16896
rect 14704 16836 14708 16892
rect 14708 16836 14764 16892
rect 14764 16836 14768 16892
rect 14704 16832 14768 16836
rect 14784 16892 14848 16896
rect 14784 16836 14788 16892
rect 14788 16836 14844 16892
rect 14844 16836 14848 16892
rect 14784 16832 14848 16836
rect 19259 16892 19323 16896
rect 19259 16836 19263 16892
rect 19263 16836 19319 16892
rect 19319 16836 19323 16892
rect 19259 16832 19323 16836
rect 19339 16892 19403 16896
rect 19339 16836 19343 16892
rect 19343 16836 19399 16892
rect 19399 16836 19403 16892
rect 19339 16832 19403 16836
rect 19419 16892 19483 16896
rect 19419 16836 19423 16892
rect 19423 16836 19479 16892
rect 19479 16836 19483 16892
rect 19419 16832 19483 16836
rect 19499 16892 19563 16896
rect 19499 16836 19503 16892
rect 19503 16836 19559 16892
rect 19559 16836 19563 16892
rect 19499 16832 19563 16836
rect 2757 16348 2821 16352
rect 2757 16292 2761 16348
rect 2761 16292 2817 16348
rect 2817 16292 2821 16348
rect 2757 16288 2821 16292
rect 2837 16348 2901 16352
rect 2837 16292 2841 16348
rect 2841 16292 2897 16348
rect 2897 16292 2901 16348
rect 2837 16288 2901 16292
rect 2917 16348 2981 16352
rect 2917 16292 2921 16348
rect 2921 16292 2977 16348
rect 2977 16292 2981 16348
rect 2917 16288 2981 16292
rect 2997 16348 3061 16352
rect 2997 16292 3001 16348
rect 3001 16292 3057 16348
rect 3057 16292 3061 16348
rect 2997 16288 3061 16292
rect 7472 16348 7536 16352
rect 7472 16292 7476 16348
rect 7476 16292 7532 16348
rect 7532 16292 7536 16348
rect 7472 16288 7536 16292
rect 7552 16348 7616 16352
rect 7552 16292 7556 16348
rect 7556 16292 7612 16348
rect 7612 16292 7616 16348
rect 7552 16288 7616 16292
rect 7632 16348 7696 16352
rect 7632 16292 7636 16348
rect 7636 16292 7692 16348
rect 7692 16292 7696 16348
rect 7632 16288 7696 16292
rect 7712 16348 7776 16352
rect 7712 16292 7716 16348
rect 7716 16292 7772 16348
rect 7772 16292 7776 16348
rect 7712 16288 7776 16292
rect 12187 16348 12251 16352
rect 12187 16292 12191 16348
rect 12191 16292 12247 16348
rect 12247 16292 12251 16348
rect 12187 16288 12251 16292
rect 12267 16348 12331 16352
rect 12267 16292 12271 16348
rect 12271 16292 12327 16348
rect 12327 16292 12331 16348
rect 12267 16288 12331 16292
rect 12347 16348 12411 16352
rect 12347 16292 12351 16348
rect 12351 16292 12407 16348
rect 12407 16292 12411 16348
rect 12347 16288 12411 16292
rect 12427 16348 12491 16352
rect 12427 16292 12431 16348
rect 12431 16292 12487 16348
rect 12487 16292 12491 16348
rect 12427 16288 12491 16292
rect 16902 16348 16966 16352
rect 16902 16292 16906 16348
rect 16906 16292 16962 16348
rect 16962 16292 16966 16348
rect 16902 16288 16966 16292
rect 16982 16348 17046 16352
rect 16982 16292 16986 16348
rect 16986 16292 17042 16348
rect 17042 16292 17046 16348
rect 16982 16288 17046 16292
rect 17062 16348 17126 16352
rect 17062 16292 17066 16348
rect 17066 16292 17122 16348
rect 17122 16292 17126 16348
rect 17062 16288 17126 16292
rect 17142 16348 17206 16352
rect 17142 16292 17146 16348
rect 17146 16292 17202 16348
rect 17202 16292 17206 16348
rect 17142 16288 17206 16292
rect 5114 15804 5178 15808
rect 5114 15748 5118 15804
rect 5118 15748 5174 15804
rect 5174 15748 5178 15804
rect 5114 15744 5178 15748
rect 5194 15804 5258 15808
rect 5194 15748 5198 15804
rect 5198 15748 5254 15804
rect 5254 15748 5258 15804
rect 5194 15744 5258 15748
rect 5274 15804 5338 15808
rect 5274 15748 5278 15804
rect 5278 15748 5334 15804
rect 5334 15748 5338 15804
rect 5274 15744 5338 15748
rect 5354 15804 5418 15808
rect 5354 15748 5358 15804
rect 5358 15748 5414 15804
rect 5414 15748 5418 15804
rect 5354 15744 5418 15748
rect 9829 15804 9893 15808
rect 9829 15748 9833 15804
rect 9833 15748 9889 15804
rect 9889 15748 9893 15804
rect 9829 15744 9893 15748
rect 9909 15804 9973 15808
rect 9909 15748 9913 15804
rect 9913 15748 9969 15804
rect 9969 15748 9973 15804
rect 9909 15744 9973 15748
rect 9989 15804 10053 15808
rect 9989 15748 9993 15804
rect 9993 15748 10049 15804
rect 10049 15748 10053 15804
rect 9989 15744 10053 15748
rect 10069 15804 10133 15808
rect 10069 15748 10073 15804
rect 10073 15748 10129 15804
rect 10129 15748 10133 15804
rect 10069 15744 10133 15748
rect 14544 15804 14608 15808
rect 14544 15748 14548 15804
rect 14548 15748 14604 15804
rect 14604 15748 14608 15804
rect 14544 15744 14608 15748
rect 14624 15804 14688 15808
rect 14624 15748 14628 15804
rect 14628 15748 14684 15804
rect 14684 15748 14688 15804
rect 14624 15744 14688 15748
rect 14704 15804 14768 15808
rect 14704 15748 14708 15804
rect 14708 15748 14764 15804
rect 14764 15748 14768 15804
rect 14704 15744 14768 15748
rect 14784 15804 14848 15808
rect 14784 15748 14788 15804
rect 14788 15748 14844 15804
rect 14844 15748 14848 15804
rect 14784 15744 14848 15748
rect 19259 15804 19323 15808
rect 19259 15748 19263 15804
rect 19263 15748 19319 15804
rect 19319 15748 19323 15804
rect 19259 15744 19323 15748
rect 19339 15804 19403 15808
rect 19339 15748 19343 15804
rect 19343 15748 19399 15804
rect 19399 15748 19403 15804
rect 19339 15744 19403 15748
rect 19419 15804 19483 15808
rect 19419 15748 19423 15804
rect 19423 15748 19479 15804
rect 19479 15748 19483 15804
rect 19419 15744 19483 15748
rect 19499 15804 19563 15808
rect 19499 15748 19503 15804
rect 19503 15748 19559 15804
rect 19559 15748 19563 15804
rect 19499 15744 19563 15748
rect 2757 15260 2821 15264
rect 2757 15204 2761 15260
rect 2761 15204 2817 15260
rect 2817 15204 2821 15260
rect 2757 15200 2821 15204
rect 2837 15260 2901 15264
rect 2837 15204 2841 15260
rect 2841 15204 2897 15260
rect 2897 15204 2901 15260
rect 2837 15200 2901 15204
rect 2917 15260 2981 15264
rect 2917 15204 2921 15260
rect 2921 15204 2977 15260
rect 2977 15204 2981 15260
rect 2917 15200 2981 15204
rect 2997 15260 3061 15264
rect 2997 15204 3001 15260
rect 3001 15204 3057 15260
rect 3057 15204 3061 15260
rect 2997 15200 3061 15204
rect 7472 15260 7536 15264
rect 7472 15204 7476 15260
rect 7476 15204 7532 15260
rect 7532 15204 7536 15260
rect 7472 15200 7536 15204
rect 7552 15260 7616 15264
rect 7552 15204 7556 15260
rect 7556 15204 7612 15260
rect 7612 15204 7616 15260
rect 7552 15200 7616 15204
rect 7632 15260 7696 15264
rect 7632 15204 7636 15260
rect 7636 15204 7692 15260
rect 7692 15204 7696 15260
rect 7632 15200 7696 15204
rect 7712 15260 7776 15264
rect 7712 15204 7716 15260
rect 7716 15204 7772 15260
rect 7772 15204 7776 15260
rect 7712 15200 7776 15204
rect 12187 15260 12251 15264
rect 12187 15204 12191 15260
rect 12191 15204 12247 15260
rect 12247 15204 12251 15260
rect 12187 15200 12251 15204
rect 12267 15260 12331 15264
rect 12267 15204 12271 15260
rect 12271 15204 12327 15260
rect 12327 15204 12331 15260
rect 12267 15200 12331 15204
rect 12347 15260 12411 15264
rect 12347 15204 12351 15260
rect 12351 15204 12407 15260
rect 12407 15204 12411 15260
rect 12347 15200 12411 15204
rect 12427 15260 12491 15264
rect 12427 15204 12431 15260
rect 12431 15204 12487 15260
rect 12487 15204 12491 15260
rect 12427 15200 12491 15204
rect 16902 15260 16966 15264
rect 16902 15204 16906 15260
rect 16906 15204 16962 15260
rect 16962 15204 16966 15260
rect 16902 15200 16966 15204
rect 16982 15260 17046 15264
rect 16982 15204 16986 15260
rect 16986 15204 17042 15260
rect 17042 15204 17046 15260
rect 16982 15200 17046 15204
rect 17062 15260 17126 15264
rect 17062 15204 17066 15260
rect 17066 15204 17122 15260
rect 17122 15204 17126 15260
rect 17062 15200 17126 15204
rect 17142 15260 17206 15264
rect 17142 15204 17146 15260
rect 17146 15204 17202 15260
rect 17202 15204 17206 15260
rect 17142 15200 17206 15204
rect 5114 14716 5178 14720
rect 5114 14660 5118 14716
rect 5118 14660 5174 14716
rect 5174 14660 5178 14716
rect 5114 14656 5178 14660
rect 5194 14716 5258 14720
rect 5194 14660 5198 14716
rect 5198 14660 5254 14716
rect 5254 14660 5258 14716
rect 5194 14656 5258 14660
rect 5274 14716 5338 14720
rect 5274 14660 5278 14716
rect 5278 14660 5334 14716
rect 5334 14660 5338 14716
rect 5274 14656 5338 14660
rect 5354 14716 5418 14720
rect 5354 14660 5358 14716
rect 5358 14660 5414 14716
rect 5414 14660 5418 14716
rect 5354 14656 5418 14660
rect 9829 14716 9893 14720
rect 9829 14660 9833 14716
rect 9833 14660 9889 14716
rect 9889 14660 9893 14716
rect 9829 14656 9893 14660
rect 9909 14716 9973 14720
rect 9909 14660 9913 14716
rect 9913 14660 9969 14716
rect 9969 14660 9973 14716
rect 9909 14656 9973 14660
rect 9989 14716 10053 14720
rect 9989 14660 9993 14716
rect 9993 14660 10049 14716
rect 10049 14660 10053 14716
rect 9989 14656 10053 14660
rect 10069 14716 10133 14720
rect 10069 14660 10073 14716
rect 10073 14660 10129 14716
rect 10129 14660 10133 14716
rect 10069 14656 10133 14660
rect 14544 14716 14608 14720
rect 14544 14660 14548 14716
rect 14548 14660 14604 14716
rect 14604 14660 14608 14716
rect 14544 14656 14608 14660
rect 14624 14716 14688 14720
rect 14624 14660 14628 14716
rect 14628 14660 14684 14716
rect 14684 14660 14688 14716
rect 14624 14656 14688 14660
rect 14704 14716 14768 14720
rect 14704 14660 14708 14716
rect 14708 14660 14764 14716
rect 14764 14660 14768 14716
rect 14704 14656 14768 14660
rect 14784 14716 14848 14720
rect 14784 14660 14788 14716
rect 14788 14660 14844 14716
rect 14844 14660 14848 14716
rect 14784 14656 14848 14660
rect 19259 14716 19323 14720
rect 19259 14660 19263 14716
rect 19263 14660 19319 14716
rect 19319 14660 19323 14716
rect 19259 14656 19323 14660
rect 19339 14716 19403 14720
rect 19339 14660 19343 14716
rect 19343 14660 19399 14716
rect 19399 14660 19403 14716
rect 19339 14656 19403 14660
rect 19419 14716 19483 14720
rect 19419 14660 19423 14716
rect 19423 14660 19479 14716
rect 19479 14660 19483 14716
rect 19419 14656 19483 14660
rect 19499 14716 19563 14720
rect 19499 14660 19503 14716
rect 19503 14660 19559 14716
rect 19559 14660 19563 14716
rect 19499 14656 19563 14660
rect 2757 14172 2821 14176
rect 2757 14116 2761 14172
rect 2761 14116 2817 14172
rect 2817 14116 2821 14172
rect 2757 14112 2821 14116
rect 2837 14172 2901 14176
rect 2837 14116 2841 14172
rect 2841 14116 2897 14172
rect 2897 14116 2901 14172
rect 2837 14112 2901 14116
rect 2917 14172 2981 14176
rect 2917 14116 2921 14172
rect 2921 14116 2977 14172
rect 2977 14116 2981 14172
rect 2917 14112 2981 14116
rect 2997 14172 3061 14176
rect 2997 14116 3001 14172
rect 3001 14116 3057 14172
rect 3057 14116 3061 14172
rect 2997 14112 3061 14116
rect 7472 14172 7536 14176
rect 7472 14116 7476 14172
rect 7476 14116 7532 14172
rect 7532 14116 7536 14172
rect 7472 14112 7536 14116
rect 7552 14172 7616 14176
rect 7552 14116 7556 14172
rect 7556 14116 7612 14172
rect 7612 14116 7616 14172
rect 7552 14112 7616 14116
rect 7632 14172 7696 14176
rect 7632 14116 7636 14172
rect 7636 14116 7692 14172
rect 7692 14116 7696 14172
rect 7632 14112 7696 14116
rect 7712 14172 7776 14176
rect 7712 14116 7716 14172
rect 7716 14116 7772 14172
rect 7772 14116 7776 14172
rect 7712 14112 7776 14116
rect 12187 14172 12251 14176
rect 12187 14116 12191 14172
rect 12191 14116 12247 14172
rect 12247 14116 12251 14172
rect 12187 14112 12251 14116
rect 12267 14172 12331 14176
rect 12267 14116 12271 14172
rect 12271 14116 12327 14172
rect 12327 14116 12331 14172
rect 12267 14112 12331 14116
rect 12347 14172 12411 14176
rect 12347 14116 12351 14172
rect 12351 14116 12407 14172
rect 12407 14116 12411 14172
rect 12347 14112 12411 14116
rect 12427 14172 12491 14176
rect 12427 14116 12431 14172
rect 12431 14116 12487 14172
rect 12487 14116 12491 14172
rect 12427 14112 12491 14116
rect 16902 14172 16966 14176
rect 16902 14116 16906 14172
rect 16906 14116 16962 14172
rect 16962 14116 16966 14172
rect 16902 14112 16966 14116
rect 16982 14172 17046 14176
rect 16982 14116 16986 14172
rect 16986 14116 17042 14172
rect 17042 14116 17046 14172
rect 16982 14112 17046 14116
rect 17062 14172 17126 14176
rect 17062 14116 17066 14172
rect 17066 14116 17122 14172
rect 17122 14116 17126 14172
rect 17062 14112 17126 14116
rect 17142 14172 17206 14176
rect 17142 14116 17146 14172
rect 17146 14116 17202 14172
rect 17202 14116 17206 14172
rect 17142 14112 17206 14116
rect 5114 13628 5178 13632
rect 5114 13572 5118 13628
rect 5118 13572 5174 13628
rect 5174 13572 5178 13628
rect 5114 13568 5178 13572
rect 5194 13628 5258 13632
rect 5194 13572 5198 13628
rect 5198 13572 5254 13628
rect 5254 13572 5258 13628
rect 5194 13568 5258 13572
rect 5274 13628 5338 13632
rect 5274 13572 5278 13628
rect 5278 13572 5334 13628
rect 5334 13572 5338 13628
rect 5274 13568 5338 13572
rect 5354 13628 5418 13632
rect 5354 13572 5358 13628
rect 5358 13572 5414 13628
rect 5414 13572 5418 13628
rect 5354 13568 5418 13572
rect 9829 13628 9893 13632
rect 9829 13572 9833 13628
rect 9833 13572 9889 13628
rect 9889 13572 9893 13628
rect 9829 13568 9893 13572
rect 9909 13628 9973 13632
rect 9909 13572 9913 13628
rect 9913 13572 9969 13628
rect 9969 13572 9973 13628
rect 9909 13568 9973 13572
rect 9989 13628 10053 13632
rect 9989 13572 9993 13628
rect 9993 13572 10049 13628
rect 10049 13572 10053 13628
rect 9989 13568 10053 13572
rect 10069 13628 10133 13632
rect 10069 13572 10073 13628
rect 10073 13572 10129 13628
rect 10129 13572 10133 13628
rect 10069 13568 10133 13572
rect 14544 13628 14608 13632
rect 14544 13572 14548 13628
rect 14548 13572 14604 13628
rect 14604 13572 14608 13628
rect 14544 13568 14608 13572
rect 14624 13628 14688 13632
rect 14624 13572 14628 13628
rect 14628 13572 14684 13628
rect 14684 13572 14688 13628
rect 14624 13568 14688 13572
rect 14704 13628 14768 13632
rect 14704 13572 14708 13628
rect 14708 13572 14764 13628
rect 14764 13572 14768 13628
rect 14704 13568 14768 13572
rect 14784 13628 14848 13632
rect 14784 13572 14788 13628
rect 14788 13572 14844 13628
rect 14844 13572 14848 13628
rect 14784 13568 14848 13572
rect 19259 13628 19323 13632
rect 19259 13572 19263 13628
rect 19263 13572 19319 13628
rect 19319 13572 19323 13628
rect 19259 13568 19323 13572
rect 19339 13628 19403 13632
rect 19339 13572 19343 13628
rect 19343 13572 19399 13628
rect 19399 13572 19403 13628
rect 19339 13568 19403 13572
rect 19419 13628 19483 13632
rect 19419 13572 19423 13628
rect 19423 13572 19479 13628
rect 19479 13572 19483 13628
rect 19419 13568 19483 13572
rect 19499 13628 19563 13632
rect 19499 13572 19503 13628
rect 19503 13572 19559 13628
rect 19559 13572 19563 13628
rect 19499 13568 19563 13572
rect 2757 13084 2821 13088
rect 2757 13028 2761 13084
rect 2761 13028 2817 13084
rect 2817 13028 2821 13084
rect 2757 13024 2821 13028
rect 2837 13084 2901 13088
rect 2837 13028 2841 13084
rect 2841 13028 2897 13084
rect 2897 13028 2901 13084
rect 2837 13024 2901 13028
rect 2917 13084 2981 13088
rect 2917 13028 2921 13084
rect 2921 13028 2977 13084
rect 2977 13028 2981 13084
rect 2917 13024 2981 13028
rect 2997 13084 3061 13088
rect 2997 13028 3001 13084
rect 3001 13028 3057 13084
rect 3057 13028 3061 13084
rect 2997 13024 3061 13028
rect 7472 13084 7536 13088
rect 7472 13028 7476 13084
rect 7476 13028 7532 13084
rect 7532 13028 7536 13084
rect 7472 13024 7536 13028
rect 7552 13084 7616 13088
rect 7552 13028 7556 13084
rect 7556 13028 7612 13084
rect 7612 13028 7616 13084
rect 7552 13024 7616 13028
rect 7632 13084 7696 13088
rect 7632 13028 7636 13084
rect 7636 13028 7692 13084
rect 7692 13028 7696 13084
rect 7632 13024 7696 13028
rect 7712 13084 7776 13088
rect 7712 13028 7716 13084
rect 7716 13028 7772 13084
rect 7772 13028 7776 13084
rect 7712 13024 7776 13028
rect 12187 13084 12251 13088
rect 12187 13028 12191 13084
rect 12191 13028 12247 13084
rect 12247 13028 12251 13084
rect 12187 13024 12251 13028
rect 12267 13084 12331 13088
rect 12267 13028 12271 13084
rect 12271 13028 12327 13084
rect 12327 13028 12331 13084
rect 12267 13024 12331 13028
rect 12347 13084 12411 13088
rect 12347 13028 12351 13084
rect 12351 13028 12407 13084
rect 12407 13028 12411 13084
rect 12347 13024 12411 13028
rect 12427 13084 12491 13088
rect 12427 13028 12431 13084
rect 12431 13028 12487 13084
rect 12487 13028 12491 13084
rect 12427 13024 12491 13028
rect 16902 13084 16966 13088
rect 16902 13028 16906 13084
rect 16906 13028 16962 13084
rect 16962 13028 16966 13084
rect 16902 13024 16966 13028
rect 16982 13084 17046 13088
rect 16982 13028 16986 13084
rect 16986 13028 17042 13084
rect 17042 13028 17046 13084
rect 16982 13024 17046 13028
rect 17062 13084 17126 13088
rect 17062 13028 17066 13084
rect 17066 13028 17122 13084
rect 17122 13028 17126 13084
rect 17062 13024 17126 13028
rect 17142 13084 17206 13088
rect 17142 13028 17146 13084
rect 17146 13028 17202 13084
rect 17202 13028 17206 13084
rect 17142 13024 17206 13028
rect 5114 12540 5178 12544
rect 5114 12484 5118 12540
rect 5118 12484 5174 12540
rect 5174 12484 5178 12540
rect 5114 12480 5178 12484
rect 5194 12540 5258 12544
rect 5194 12484 5198 12540
rect 5198 12484 5254 12540
rect 5254 12484 5258 12540
rect 5194 12480 5258 12484
rect 5274 12540 5338 12544
rect 5274 12484 5278 12540
rect 5278 12484 5334 12540
rect 5334 12484 5338 12540
rect 5274 12480 5338 12484
rect 5354 12540 5418 12544
rect 5354 12484 5358 12540
rect 5358 12484 5414 12540
rect 5414 12484 5418 12540
rect 5354 12480 5418 12484
rect 9829 12540 9893 12544
rect 9829 12484 9833 12540
rect 9833 12484 9889 12540
rect 9889 12484 9893 12540
rect 9829 12480 9893 12484
rect 9909 12540 9973 12544
rect 9909 12484 9913 12540
rect 9913 12484 9969 12540
rect 9969 12484 9973 12540
rect 9909 12480 9973 12484
rect 9989 12540 10053 12544
rect 9989 12484 9993 12540
rect 9993 12484 10049 12540
rect 10049 12484 10053 12540
rect 9989 12480 10053 12484
rect 10069 12540 10133 12544
rect 10069 12484 10073 12540
rect 10073 12484 10129 12540
rect 10129 12484 10133 12540
rect 10069 12480 10133 12484
rect 14544 12540 14608 12544
rect 14544 12484 14548 12540
rect 14548 12484 14604 12540
rect 14604 12484 14608 12540
rect 14544 12480 14608 12484
rect 14624 12540 14688 12544
rect 14624 12484 14628 12540
rect 14628 12484 14684 12540
rect 14684 12484 14688 12540
rect 14624 12480 14688 12484
rect 14704 12540 14768 12544
rect 14704 12484 14708 12540
rect 14708 12484 14764 12540
rect 14764 12484 14768 12540
rect 14704 12480 14768 12484
rect 14784 12540 14848 12544
rect 14784 12484 14788 12540
rect 14788 12484 14844 12540
rect 14844 12484 14848 12540
rect 14784 12480 14848 12484
rect 19259 12540 19323 12544
rect 19259 12484 19263 12540
rect 19263 12484 19319 12540
rect 19319 12484 19323 12540
rect 19259 12480 19323 12484
rect 19339 12540 19403 12544
rect 19339 12484 19343 12540
rect 19343 12484 19399 12540
rect 19399 12484 19403 12540
rect 19339 12480 19403 12484
rect 19419 12540 19483 12544
rect 19419 12484 19423 12540
rect 19423 12484 19479 12540
rect 19479 12484 19483 12540
rect 19419 12480 19483 12484
rect 19499 12540 19563 12544
rect 19499 12484 19503 12540
rect 19503 12484 19559 12540
rect 19559 12484 19563 12540
rect 19499 12480 19563 12484
rect 2757 11996 2821 12000
rect 2757 11940 2761 11996
rect 2761 11940 2817 11996
rect 2817 11940 2821 11996
rect 2757 11936 2821 11940
rect 2837 11996 2901 12000
rect 2837 11940 2841 11996
rect 2841 11940 2897 11996
rect 2897 11940 2901 11996
rect 2837 11936 2901 11940
rect 2917 11996 2981 12000
rect 2917 11940 2921 11996
rect 2921 11940 2977 11996
rect 2977 11940 2981 11996
rect 2917 11936 2981 11940
rect 2997 11996 3061 12000
rect 2997 11940 3001 11996
rect 3001 11940 3057 11996
rect 3057 11940 3061 11996
rect 2997 11936 3061 11940
rect 7472 11996 7536 12000
rect 7472 11940 7476 11996
rect 7476 11940 7532 11996
rect 7532 11940 7536 11996
rect 7472 11936 7536 11940
rect 7552 11996 7616 12000
rect 7552 11940 7556 11996
rect 7556 11940 7612 11996
rect 7612 11940 7616 11996
rect 7552 11936 7616 11940
rect 7632 11996 7696 12000
rect 7632 11940 7636 11996
rect 7636 11940 7692 11996
rect 7692 11940 7696 11996
rect 7632 11936 7696 11940
rect 7712 11996 7776 12000
rect 7712 11940 7716 11996
rect 7716 11940 7772 11996
rect 7772 11940 7776 11996
rect 7712 11936 7776 11940
rect 12187 11996 12251 12000
rect 12187 11940 12191 11996
rect 12191 11940 12247 11996
rect 12247 11940 12251 11996
rect 12187 11936 12251 11940
rect 12267 11996 12331 12000
rect 12267 11940 12271 11996
rect 12271 11940 12327 11996
rect 12327 11940 12331 11996
rect 12267 11936 12331 11940
rect 12347 11996 12411 12000
rect 12347 11940 12351 11996
rect 12351 11940 12407 11996
rect 12407 11940 12411 11996
rect 12347 11936 12411 11940
rect 12427 11996 12491 12000
rect 12427 11940 12431 11996
rect 12431 11940 12487 11996
rect 12487 11940 12491 11996
rect 12427 11936 12491 11940
rect 16902 11996 16966 12000
rect 16902 11940 16906 11996
rect 16906 11940 16962 11996
rect 16962 11940 16966 11996
rect 16902 11936 16966 11940
rect 16982 11996 17046 12000
rect 16982 11940 16986 11996
rect 16986 11940 17042 11996
rect 17042 11940 17046 11996
rect 16982 11936 17046 11940
rect 17062 11996 17126 12000
rect 17062 11940 17066 11996
rect 17066 11940 17122 11996
rect 17122 11940 17126 11996
rect 17062 11936 17126 11940
rect 17142 11996 17206 12000
rect 17142 11940 17146 11996
rect 17146 11940 17202 11996
rect 17202 11940 17206 11996
rect 17142 11936 17206 11940
rect 5114 11452 5178 11456
rect 5114 11396 5118 11452
rect 5118 11396 5174 11452
rect 5174 11396 5178 11452
rect 5114 11392 5178 11396
rect 5194 11452 5258 11456
rect 5194 11396 5198 11452
rect 5198 11396 5254 11452
rect 5254 11396 5258 11452
rect 5194 11392 5258 11396
rect 5274 11452 5338 11456
rect 5274 11396 5278 11452
rect 5278 11396 5334 11452
rect 5334 11396 5338 11452
rect 5274 11392 5338 11396
rect 5354 11452 5418 11456
rect 5354 11396 5358 11452
rect 5358 11396 5414 11452
rect 5414 11396 5418 11452
rect 5354 11392 5418 11396
rect 9829 11452 9893 11456
rect 9829 11396 9833 11452
rect 9833 11396 9889 11452
rect 9889 11396 9893 11452
rect 9829 11392 9893 11396
rect 9909 11452 9973 11456
rect 9909 11396 9913 11452
rect 9913 11396 9969 11452
rect 9969 11396 9973 11452
rect 9909 11392 9973 11396
rect 9989 11452 10053 11456
rect 9989 11396 9993 11452
rect 9993 11396 10049 11452
rect 10049 11396 10053 11452
rect 9989 11392 10053 11396
rect 10069 11452 10133 11456
rect 10069 11396 10073 11452
rect 10073 11396 10129 11452
rect 10129 11396 10133 11452
rect 10069 11392 10133 11396
rect 14544 11452 14608 11456
rect 14544 11396 14548 11452
rect 14548 11396 14604 11452
rect 14604 11396 14608 11452
rect 14544 11392 14608 11396
rect 14624 11452 14688 11456
rect 14624 11396 14628 11452
rect 14628 11396 14684 11452
rect 14684 11396 14688 11452
rect 14624 11392 14688 11396
rect 14704 11452 14768 11456
rect 14704 11396 14708 11452
rect 14708 11396 14764 11452
rect 14764 11396 14768 11452
rect 14704 11392 14768 11396
rect 14784 11452 14848 11456
rect 14784 11396 14788 11452
rect 14788 11396 14844 11452
rect 14844 11396 14848 11452
rect 14784 11392 14848 11396
rect 19259 11452 19323 11456
rect 19259 11396 19263 11452
rect 19263 11396 19319 11452
rect 19319 11396 19323 11452
rect 19259 11392 19323 11396
rect 19339 11452 19403 11456
rect 19339 11396 19343 11452
rect 19343 11396 19399 11452
rect 19399 11396 19403 11452
rect 19339 11392 19403 11396
rect 19419 11452 19483 11456
rect 19419 11396 19423 11452
rect 19423 11396 19479 11452
rect 19479 11396 19483 11452
rect 19419 11392 19483 11396
rect 19499 11452 19563 11456
rect 19499 11396 19503 11452
rect 19503 11396 19559 11452
rect 19559 11396 19563 11452
rect 19499 11392 19563 11396
rect 2757 10908 2821 10912
rect 2757 10852 2761 10908
rect 2761 10852 2817 10908
rect 2817 10852 2821 10908
rect 2757 10848 2821 10852
rect 2837 10908 2901 10912
rect 2837 10852 2841 10908
rect 2841 10852 2897 10908
rect 2897 10852 2901 10908
rect 2837 10848 2901 10852
rect 2917 10908 2981 10912
rect 2917 10852 2921 10908
rect 2921 10852 2977 10908
rect 2977 10852 2981 10908
rect 2917 10848 2981 10852
rect 2997 10908 3061 10912
rect 2997 10852 3001 10908
rect 3001 10852 3057 10908
rect 3057 10852 3061 10908
rect 2997 10848 3061 10852
rect 7472 10908 7536 10912
rect 7472 10852 7476 10908
rect 7476 10852 7532 10908
rect 7532 10852 7536 10908
rect 7472 10848 7536 10852
rect 7552 10908 7616 10912
rect 7552 10852 7556 10908
rect 7556 10852 7612 10908
rect 7612 10852 7616 10908
rect 7552 10848 7616 10852
rect 7632 10908 7696 10912
rect 7632 10852 7636 10908
rect 7636 10852 7692 10908
rect 7692 10852 7696 10908
rect 7632 10848 7696 10852
rect 7712 10908 7776 10912
rect 7712 10852 7716 10908
rect 7716 10852 7772 10908
rect 7772 10852 7776 10908
rect 7712 10848 7776 10852
rect 12187 10908 12251 10912
rect 12187 10852 12191 10908
rect 12191 10852 12247 10908
rect 12247 10852 12251 10908
rect 12187 10848 12251 10852
rect 12267 10908 12331 10912
rect 12267 10852 12271 10908
rect 12271 10852 12327 10908
rect 12327 10852 12331 10908
rect 12267 10848 12331 10852
rect 12347 10908 12411 10912
rect 12347 10852 12351 10908
rect 12351 10852 12407 10908
rect 12407 10852 12411 10908
rect 12347 10848 12411 10852
rect 12427 10908 12491 10912
rect 12427 10852 12431 10908
rect 12431 10852 12487 10908
rect 12487 10852 12491 10908
rect 12427 10848 12491 10852
rect 16902 10908 16966 10912
rect 16902 10852 16906 10908
rect 16906 10852 16962 10908
rect 16962 10852 16966 10908
rect 16902 10848 16966 10852
rect 16982 10908 17046 10912
rect 16982 10852 16986 10908
rect 16986 10852 17042 10908
rect 17042 10852 17046 10908
rect 16982 10848 17046 10852
rect 17062 10908 17126 10912
rect 17062 10852 17066 10908
rect 17066 10852 17122 10908
rect 17122 10852 17126 10908
rect 17062 10848 17126 10852
rect 17142 10908 17206 10912
rect 17142 10852 17146 10908
rect 17146 10852 17202 10908
rect 17202 10852 17206 10908
rect 17142 10848 17206 10852
rect 5114 10364 5178 10368
rect 5114 10308 5118 10364
rect 5118 10308 5174 10364
rect 5174 10308 5178 10364
rect 5114 10304 5178 10308
rect 5194 10364 5258 10368
rect 5194 10308 5198 10364
rect 5198 10308 5254 10364
rect 5254 10308 5258 10364
rect 5194 10304 5258 10308
rect 5274 10364 5338 10368
rect 5274 10308 5278 10364
rect 5278 10308 5334 10364
rect 5334 10308 5338 10364
rect 5274 10304 5338 10308
rect 5354 10364 5418 10368
rect 5354 10308 5358 10364
rect 5358 10308 5414 10364
rect 5414 10308 5418 10364
rect 5354 10304 5418 10308
rect 9829 10364 9893 10368
rect 9829 10308 9833 10364
rect 9833 10308 9889 10364
rect 9889 10308 9893 10364
rect 9829 10304 9893 10308
rect 9909 10364 9973 10368
rect 9909 10308 9913 10364
rect 9913 10308 9969 10364
rect 9969 10308 9973 10364
rect 9909 10304 9973 10308
rect 9989 10364 10053 10368
rect 9989 10308 9993 10364
rect 9993 10308 10049 10364
rect 10049 10308 10053 10364
rect 9989 10304 10053 10308
rect 10069 10364 10133 10368
rect 10069 10308 10073 10364
rect 10073 10308 10129 10364
rect 10129 10308 10133 10364
rect 10069 10304 10133 10308
rect 14544 10364 14608 10368
rect 14544 10308 14548 10364
rect 14548 10308 14604 10364
rect 14604 10308 14608 10364
rect 14544 10304 14608 10308
rect 14624 10364 14688 10368
rect 14624 10308 14628 10364
rect 14628 10308 14684 10364
rect 14684 10308 14688 10364
rect 14624 10304 14688 10308
rect 14704 10364 14768 10368
rect 14704 10308 14708 10364
rect 14708 10308 14764 10364
rect 14764 10308 14768 10364
rect 14704 10304 14768 10308
rect 14784 10364 14848 10368
rect 14784 10308 14788 10364
rect 14788 10308 14844 10364
rect 14844 10308 14848 10364
rect 14784 10304 14848 10308
rect 19259 10364 19323 10368
rect 19259 10308 19263 10364
rect 19263 10308 19319 10364
rect 19319 10308 19323 10364
rect 19259 10304 19323 10308
rect 19339 10364 19403 10368
rect 19339 10308 19343 10364
rect 19343 10308 19399 10364
rect 19399 10308 19403 10364
rect 19339 10304 19403 10308
rect 19419 10364 19483 10368
rect 19419 10308 19423 10364
rect 19423 10308 19479 10364
rect 19479 10308 19483 10364
rect 19419 10304 19483 10308
rect 19499 10364 19563 10368
rect 19499 10308 19503 10364
rect 19503 10308 19559 10364
rect 19559 10308 19563 10364
rect 19499 10304 19563 10308
rect 2757 9820 2821 9824
rect 2757 9764 2761 9820
rect 2761 9764 2817 9820
rect 2817 9764 2821 9820
rect 2757 9760 2821 9764
rect 2837 9820 2901 9824
rect 2837 9764 2841 9820
rect 2841 9764 2897 9820
rect 2897 9764 2901 9820
rect 2837 9760 2901 9764
rect 2917 9820 2981 9824
rect 2917 9764 2921 9820
rect 2921 9764 2977 9820
rect 2977 9764 2981 9820
rect 2917 9760 2981 9764
rect 2997 9820 3061 9824
rect 2997 9764 3001 9820
rect 3001 9764 3057 9820
rect 3057 9764 3061 9820
rect 2997 9760 3061 9764
rect 7472 9820 7536 9824
rect 7472 9764 7476 9820
rect 7476 9764 7532 9820
rect 7532 9764 7536 9820
rect 7472 9760 7536 9764
rect 7552 9820 7616 9824
rect 7552 9764 7556 9820
rect 7556 9764 7612 9820
rect 7612 9764 7616 9820
rect 7552 9760 7616 9764
rect 7632 9820 7696 9824
rect 7632 9764 7636 9820
rect 7636 9764 7692 9820
rect 7692 9764 7696 9820
rect 7632 9760 7696 9764
rect 7712 9820 7776 9824
rect 7712 9764 7716 9820
rect 7716 9764 7772 9820
rect 7772 9764 7776 9820
rect 7712 9760 7776 9764
rect 12187 9820 12251 9824
rect 12187 9764 12191 9820
rect 12191 9764 12247 9820
rect 12247 9764 12251 9820
rect 12187 9760 12251 9764
rect 12267 9820 12331 9824
rect 12267 9764 12271 9820
rect 12271 9764 12327 9820
rect 12327 9764 12331 9820
rect 12267 9760 12331 9764
rect 12347 9820 12411 9824
rect 12347 9764 12351 9820
rect 12351 9764 12407 9820
rect 12407 9764 12411 9820
rect 12347 9760 12411 9764
rect 12427 9820 12491 9824
rect 12427 9764 12431 9820
rect 12431 9764 12487 9820
rect 12487 9764 12491 9820
rect 12427 9760 12491 9764
rect 16902 9820 16966 9824
rect 16902 9764 16906 9820
rect 16906 9764 16962 9820
rect 16962 9764 16966 9820
rect 16902 9760 16966 9764
rect 16982 9820 17046 9824
rect 16982 9764 16986 9820
rect 16986 9764 17042 9820
rect 17042 9764 17046 9820
rect 16982 9760 17046 9764
rect 17062 9820 17126 9824
rect 17062 9764 17066 9820
rect 17066 9764 17122 9820
rect 17122 9764 17126 9820
rect 17062 9760 17126 9764
rect 17142 9820 17206 9824
rect 17142 9764 17146 9820
rect 17146 9764 17202 9820
rect 17202 9764 17206 9820
rect 17142 9760 17206 9764
rect 5114 9276 5178 9280
rect 5114 9220 5118 9276
rect 5118 9220 5174 9276
rect 5174 9220 5178 9276
rect 5114 9216 5178 9220
rect 5194 9276 5258 9280
rect 5194 9220 5198 9276
rect 5198 9220 5254 9276
rect 5254 9220 5258 9276
rect 5194 9216 5258 9220
rect 5274 9276 5338 9280
rect 5274 9220 5278 9276
rect 5278 9220 5334 9276
rect 5334 9220 5338 9276
rect 5274 9216 5338 9220
rect 5354 9276 5418 9280
rect 5354 9220 5358 9276
rect 5358 9220 5414 9276
rect 5414 9220 5418 9276
rect 5354 9216 5418 9220
rect 9829 9276 9893 9280
rect 9829 9220 9833 9276
rect 9833 9220 9889 9276
rect 9889 9220 9893 9276
rect 9829 9216 9893 9220
rect 9909 9276 9973 9280
rect 9909 9220 9913 9276
rect 9913 9220 9969 9276
rect 9969 9220 9973 9276
rect 9909 9216 9973 9220
rect 9989 9276 10053 9280
rect 9989 9220 9993 9276
rect 9993 9220 10049 9276
rect 10049 9220 10053 9276
rect 9989 9216 10053 9220
rect 10069 9276 10133 9280
rect 10069 9220 10073 9276
rect 10073 9220 10129 9276
rect 10129 9220 10133 9276
rect 10069 9216 10133 9220
rect 14544 9276 14608 9280
rect 14544 9220 14548 9276
rect 14548 9220 14604 9276
rect 14604 9220 14608 9276
rect 14544 9216 14608 9220
rect 14624 9276 14688 9280
rect 14624 9220 14628 9276
rect 14628 9220 14684 9276
rect 14684 9220 14688 9276
rect 14624 9216 14688 9220
rect 14704 9276 14768 9280
rect 14704 9220 14708 9276
rect 14708 9220 14764 9276
rect 14764 9220 14768 9276
rect 14704 9216 14768 9220
rect 14784 9276 14848 9280
rect 14784 9220 14788 9276
rect 14788 9220 14844 9276
rect 14844 9220 14848 9276
rect 14784 9216 14848 9220
rect 19259 9276 19323 9280
rect 19259 9220 19263 9276
rect 19263 9220 19319 9276
rect 19319 9220 19323 9276
rect 19259 9216 19323 9220
rect 19339 9276 19403 9280
rect 19339 9220 19343 9276
rect 19343 9220 19399 9276
rect 19399 9220 19403 9276
rect 19339 9216 19403 9220
rect 19419 9276 19483 9280
rect 19419 9220 19423 9276
rect 19423 9220 19479 9276
rect 19479 9220 19483 9276
rect 19419 9216 19483 9220
rect 19499 9276 19563 9280
rect 19499 9220 19503 9276
rect 19503 9220 19559 9276
rect 19559 9220 19563 9276
rect 19499 9216 19563 9220
rect 2757 8732 2821 8736
rect 2757 8676 2761 8732
rect 2761 8676 2817 8732
rect 2817 8676 2821 8732
rect 2757 8672 2821 8676
rect 2837 8732 2901 8736
rect 2837 8676 2841 8732
rect 2841 8676 2897 8732
rect 2897 8676 2901 8732
rect 2837 8672 2901 8676
rect 2917 8732 2981 8736
rect 2917 8676 2921 8732
rect 2921 8676 2977 8732
rect 2977 8676 2981 8732
rect 2917 8672 2981 8676
rect 2997 8732 3061 8736
rect 2997 8676 3001 8732
rect 3001 8676 3057 8732
rect 3057 8676 3061 8732
rect 2997 8672 3061 8676
rect 7472 8732 7536 8736
rect 7472 8676 7476 8732
rect 7476 8676 7532 8732
rect 7532 8676 7536 8732
rect 7472 8672 7536 8676
rect 7552 8732 7616 8736
rect 7552 8676 7556 8732
rect 7556 8676 7612 8732
rect 7612 8676 7616 8732
rect 7552 8672 7616 8676
rect 7632 8732 7696 8736
rect 7632 8676 7636 8732
rect 7636 8676 7692 8732
rect 7692 8676 7696 8732
rect 7632 8672 7696 8676
rect 7712 8732 7776 8736
rect 7712 8676 7716 8732
rect 7716 8676 7772 8732
rect 7772 8676 7776 8732
rect 7712 8672 7776 8676
rect 12187 8732 12251 8736
rect 12187 8676 12191 8732
rect 12191 8676 12247 8732
rect 12247 8676 12251 8732
rect 12187 8672 12251 8676
rect 12267 8732 12331 8736
rect 12267 8676 12271 8732
rect 12271 8676 12327 8732
rect 12327 8676 12331 8732
rect 12267 8672 12331 8676
rect 12347 8732 12411 8736
rect 12347 8676 12351 8732
rect 12351 8676 12407 8732
rect 12407 8676 12411 8732
rect 12347 8672 12411 8676
rect 12427 8732 12491 8736
rect 12427 8676 12431 8732
rect 12431 8676 12487 8732
rect 12487 8676 12491 8732
rect 12427 8672 12491 8676
rect 16902 8732 16966 8736
rect 16902 8676 16906 8732
rect 16906 8676 16962 8732
rect 16962 8676 16966 8732
rect 16902 8672 16966 8676
rect 16982 8732 17046 8736
rect 16982 8676 16986 8732
rect 16986 8676 17042 8732
rect 17042 8676 17046 8732
rect 16982 8672 17046 8676
rect 17062 8732 17126 8736
rect 17062 8676 17066 8732
rect 17066 8676 17122 8732
rect 17122 8676 17126 8732
rect 17062 8672 17126 8676
rect 17142 8732 17206 8736
rect 17142 8676 17146 8732
rect 17146 8676 17202 8732
rect 17202 8676 17206 8732
rect 17142 8672 17206 8676
rect 5114 8188 5178 8192
rect 5114 8132 5118 8188
rect 5118 8132 5174 8188
rect 5174 8132 5178 8188
rect 5114 8128 5178 8132
rect 5194 8188 5258 8192
rect 5194 8132 5198 8188
rect 5198 8132 5254 8188
rect 5254 8132 5258 8188
rect 5194 8128 5258 8132
rect 5274 8188 5338 8192
rect 5274 8132 5278 8188
rect 5278 8132 5334 8188
rect 5334 8132 5338 8188
rect 5274 8128 5338 8132
rect 5354 8188 5418 8192
rect 5354 8132 5358 8188
rect 5358 8132 5414 8188
rect 5414 8132 5418 8188
rect 5354 8128 5418 8132
rect 9829 8188 9893 8192
rect 9829 8132 9833 8188
rect 9833 8132 9889 8188
rect 9889 8132 9893 8188
rect 9829 8128 9893 8132
rect 9909 8188 9973 8192
rect 9909 8132 9913 8188
rect 9913 8132 9969 8188
rect 9969 8132 9973 8188
rect 9909 8128 9973 8132
rect 9989 8188 10053 8192
rect 9989 8132 9993 8188
rect 9993 8132 10049 8188
rect 10049 8132 10053 8188
rect 9989 8128 10053 8132
rect 10069 8188 10133 8192
rect 10069 8132 10073 8188
rect 10073 8132 10129 8188
rect 10129 8132 10133 8188
rect 10069 8128 10133 8132
rect 14544 8188 14608 8192
rect 14544 8132 14548 8188
rect 14548 8132 14604 8188
rect 14604 8132 14608 8188
rect 14544 8128 14608 8132
rect 14624 8188 14688 8192
rect 14624 8132 14628 8188
rect 14628 8132 14684 8188
rect 14684 8132 14688 8188
rect 14624 8128 14688 8132
rect 14704 8188 14768 8192
rect 14704 8132 14708 8188
rect 14708 8132 14764 8188
rect 14764 8132 14768 8188
rect 14704 8128 14768 8132
rect 14784 8188 14848 8192
rect 14784 8132 14788 8188
rect 14788 8132 14844 8188
rect 14844 8132 14848 8188
rect 14784 8128 14848 8132
rect 19259 8188 19323 8192
rect 19259 8132 19263 8188
rect 19263 8132 19319 8188
rect 19319 8132 19323 8188
rect 19259 8128 19323 8132
rect 19339 8188 19403 8192
rect 19339 8132 19343 8188
rect 19343 8132 19399 8188
rect 19399 8132 19403 8188
rect 19339 8128 19403 8132
rect 19419 8188 19483 8192
rect 19419 8132 19423 8188
rect 19423 8132 19479 8188
rect 19479 8132 19483 8188
rect 19419 8128 19483 8132
rect 19499 8188 19563 8192
rect 19499 8132 19503 8188
rect 19503 8132 19559 8188
rect 19559 8132 19563 8188
rect 19499 8128 19563 8132
rect 2757 7644 2821 7648
rect 2757 7588 2761 7644
rect 2761 7588 2817 7644
rect 2817 7588 2821 7644
rect 2757 7584 2821 7588
rect 2837 7644 2901 7648
rect 2837 7588 2841 7644
rect 2841 7588 2897 7644
rect 2897 7588 2901 7644
rect 2837 7584 2901 7588
rect 2917 7644 2981 7648
rect 2917 7588 2921 7644
rect 2921 7588 2977 7644
rect 2977 7588 2981 7644
rect 2917 7584 2981 7588
rect 2997 7644 3061 7648
rect 2997 7588 3001 7644
rect 3001 7588 3057 7644
rect 3057 7588 3061 7644
rect 2997 7584 3061 7588
rect 7472 7644 7536 7648
rect 7472 7588 7476 7644
rect 7476 7588 7532 7644
rect 7532 7588 7536 7644
rect 7472 7584 7536 7588
rect 7552 7644 7616 7648
rect 7552 7588 7556 7644
rect 7556 7588 7612 7644
rect 7612 7588 7616 7644
rect 7552 7584 7616 7588
rect 7632 7644 7696 7648
rect 7632 7588 7636 7644
rect 7636 7588 7692 7644
rect 7692 7588 7696 7644
rect 7632 7584 7696 7588
rect 7712 7644 7776 7648
rect 7712 7588 7716 7644
rect 7716 7588 7772 7644
rect 7772 7588 7776 7644
rect 7712 7584 7776 7588
rect 12187 7644 12251 7648
rect 12187 7588 12191 7644
rect 12191 7588 12247 7644
rect 12247 7588 12251 7644
rect 12187 7584 12251 7588
rect 12267 7644 12331 7648
rect 12267 7588 12271 7644
rect 12271 7588 12327 7644
rect 12327 7588 12331 7644
rect 12267 7584 12331 7588
rect 12347 7644 12411 7648
rect 12347 7588 12351 7644
rect 12351 7588 12407 7644
rect 12407 7588 12411 7644
rect 12347 7584 12411 7588
rect 12427 7644 12491 7648
rect 12427 7588 12431 7644
rect 12431 7588 12487 7644
rect 12487 7588 12491 7644
rect 12427 7584 12491 7588
rect 16902 7644 16966 7648
rect 16902 7588 16906 7644
rect 16906 7588 16962 7644
rect 16962 7588 16966 7644
rect 16902 7584 16966 7588
rect 16982 7644 17046 7648
rect 16982 7588 16986 7644
rect 16986 7588 17042 7644
rect 17042 7588 17046 7644
rect 16982 7584 17046 7588
rect 17062 7644 17126 7648
rect 17062 7588 17066 7644
rect 17066 7588 17122 7644
rect 17122 7588 17126 7644
rect 17062 7584 17126 7588
rect 17142 7644 17206 7648
rect 17142 7588 17146 7644
rect 17146 7588 17202 7644
rect 17202 7588 17206 7644
rect 17142 7584 17206 7588
rect 5114 7100 5178 7104
rect 5114 7044 5118 7100
rect 5118 7044 5174 7100
rect 5174 7044 5178 7100
rect 5114 7040 5178 7044
rect 5194 7100 5258 7104
rect 5194 7044 5198 7100
rect 5198 7044 5254 7100
rect 5254 7044 5258 7100
rect 5194 7040 5258 7044
rect 5274 7100 5338 7104
rect 5274 7044 5278 7100
rect 5278 7044 5334 7100
rect 5334 7044 5338 7100
rect 5274 7040 5338 7044
rect 5354 7100 5418 7104
rect 5354 7044 5358 7100
rect 5358 7044 5414 7100
rect 5414 7044 5418 7100
rect 5354 7040 5418 7044
rect 9829 7100 9893 7104
rect 9829 7044 9833 7100
rect 9833 7044 9889 7100
rect 9889 7044 9893 7100
rect 9829 7040 9893 7044
rect 9909 7100 9973 7104
rect 9909 7044 9913 7100
rect 9913 7044 9969 7100
rect 9969 7044 9973 7100
rect 9909 7040 9973 7044
rect 9989 7100 10053 7104
rect 9989 7044 9993 7100
rect 9993 7044 10049 7100
rect 10049 7044 10053 7100
rect 9989 7040 10053 7044
rect 10069 7100 10133 7104
rect 10069 7044 10073 7100
rect 10073 7044 10129 7100
rect 10129 7044 10133 7100
rect 10069 7040 10133 7044
rect 14544 7100 14608 7104
rect 14544 7044 14548 7100
rect 14548 7044 14604 7100
rect 14604 7044 14608 7100
rect 14544 7040 14608 7044
rect 14624 7100 14688 7104
rect 14624 7044 14628 7100
rect 14628 7044 14684 7100
rect 14684 7044 14688 7100
rect 14624 7040 14688 7044
rect 14704 7100 14768 7104
rect 14704 7044 14708 7100
rect 14708 7044 14764 7100
rect 14764 7044 14768 7100
rect 14704 7040 14768 7044
rect 14784 7100 14848 7104
rect 14784 7044 14788 7100
rect 14788 7044 14844 7100
rect 14844 7044 14848 7100
rect 14784 7040 14848 7044
rect 19259 7100 19323 7104
rect 19259 7044 19263 7100
rect 19263 7044 19319 7100
rect 19319 7044 19323 7100
rect 19259 7040 19323 7044
rect 19339 7100 19403 7104
rect 19339 7044 19343 7100
rect 19343 7044 19399 7100
rect 19399 7044 19403 7100
rect 19339 7040 19403 7044
rect 19419 7100 19483 7104
rect 19419 7044 19423 7100
rect 19423 7044 19479 7100
rect 19479 7044 19483 7100
rect 19419 7040 19483 7044
rect 19499 7100 19563 7104
rect 19499 7044 19503 7100
rect 19503 7044 19559 7100
rect 19559 7044 19563 7100
rect 19499 7040 19563 7044
rect 2757 6556 2821 6560
rect 2757 6500 2761 6556
rect 2761 6500 2817 6556
rect 2817 6500 2821 6556
rect 2757 6496 2821 6500
rect 2837 6556 2901 6560
rect 2837 6500 2841 6556
rect 2841 6500 2897 6556
rect 2897 6500 2901 6556
rect 2837 6496 2901 6500
rect 2917 6556 2981 6560
rect 2917 6500 2921 6556
rect 2921 6500 2977 6556
rect 2977 6500 2981 6556
rect 2917 6496 2981 6500
rect 2997 6556 3061 6560
rect 2997 6500 3001 6556
rect 3001 6500 3057 6556
rect 3057 6500 3061 6556
rect 2997 6496 3061 6500
rect 7472 6556 7536 6560
rect 7472 6500 7476 6556
rect 7476 6500 7532 6556
rect 7532 6500 7536 6556
rect 7472 6496 7536 6500
rect 7552 6556 7616 6560
rect 7552 6500 7556 6556
rect 7556 6500 7612 6556
rect 7612 6500 7616 6556
rect 7552 6496 7616 6500
rect 7632 6556 7696 6560
rect 7632 6500 7636 6556
rect 7636 6500 7692 6556
rect 7692 6500 7696 6556
rect 7632 6496 7696 6500
rect 7712 6556 7776 6560
rect 7712 6500 7716 6556
rect 7716 6500 7772 6556
rect 7772 6500 7776 6556
rect 7712 6496 7776 6500
rect 12187 6556 12251 6560
rect 12187 6500 12191 6556
rect 12191 6500 12247 6556
rect 12247 6500 12251 6556
rect 12187 6496 12251 6500
rect 12267 6556 12331 6560
rect 12267 6500 12271 6556
rect 12271 6500 12327 6556
rect 12327 6500 12331 6556
rect 12267 6496 12331 6500
rect 12347 6556 12411 6560
rect 12347 6500 12351 6556
rect 12351 6500 12407 6556
rect 12407 6500 12411 6556
rect 12347 6496 12411 6500
rect 12427 6556 12491 6560
rect 12427 6500 12431 6556
rect 12431 6500 12487 6556
rect 12487 6500 12491 6556
rect 12427 6496 12491 6500
rect 16902 6556 16966 6560
rect 16902 6500 16906 6556
rect 16906 6500 16962 6556
rect 16962 6500 16966 6556
rect 16902 6496 16966 6500
rect 16982 6556 17046 6560
rect 16982 6500 16986 6556
rect 16986 6500 17042 6556
rect 17042 6500 17046 6556
rect 16982 6496 17046 6500
rect 17062 6556 17126 6560
rect 17062 6500 17066 6556
rect 17066 6500 17122 6556
rect 17122 6500 17126 6556
rect 17062 6496 17126 6500
rect 17142 6556 17206 6560
rect 17142 6500 17146 6556
rect 17146 6500 17202 6556
rect 17202 6500 17206 6556
rect 17142 6496 17206 6500
rect 5114 6012 5178 6016
rect 5114 5956 5118 6012
rect 5118 5956 5174 6012
rect 5174 5956 5178 6012
rect 5114 5952 5178 5956
rect 5194 6012 5258 6016
rect 5194 5956 5198 6012
rect 5198 5956 5254 6012
rect 5254 5956 5258 6012
rect 5194 5952 5258 5956
rect 5274 6012 5338 6016
rect 5274 5956 5278 6012
rect 5278 5956 5334 6012
rect 5334 5956 5338 6012
rect 5274 5952 5338 5956
rect 5354 6012 5418 6016
rect 5354 5956 5358 6012
rect 5358 5956 5414 6012
rect 5414 5956 5418 6012
rect 5354 5952 5418 5956
rect 9829 6012 9893 6016
rect 9829 5956 9833 6012
rect 9833 5956 9889 6012
rect 9889 5956 9893 6012
rect 9829 5952 9893 5956
rect 9909 6012 9973 6016
rect 9909 5956 9913 6012
rect 9913 5956 9969 6012
rect 9969 5956 9973 6012
rect 9909 5952 9973 5956
rect 9989 6012 10053 6016
rect 9989 5956 9993 6012
rect 9993 5956 10049 6012
rect 10049 5956 10053 6012
rect 9989 5952 10053 5956
rect 10069 6012 10133 6016
rect 10069 5956 10073 6012
rect 10073 5956 10129 6012
rect 10129 5956 10133 6012
rect 10069 5952 10133 5956
rect 14544 6012 14608 6016
rect 14544 5956 14548 6012
rect 14548 5956 14604 6012
rect 14604 5956 14608 6012
rect 14544 5952 14608 5956
rect 14624 6012 14688 6016
rect 14624 5956 14628 6012
rect 14628 5956 14684 6012
rect 14684 5956 14688 6012
rect 14624 5952 14688 5956
rect 14704 6012 14768 6016
rect 14704 5956 14708 6012
rect 14708 5956 14764 6012
rect 14764 5956 14768 6012
rect 14704 5952 14768 5956
rect 14784 6012 14848 6016
rect 14784 5956 14788 6012
rect 14788 5956 14844 6012
rect 14844 5956 14848 6012
rect 14784 5952 14848 5956
rect 19259 6012 19323 6016
rect 19259 5956 19263 6012
rect 19263 5956 19319 6012
rect 19319 5956 19323 6012
rect 19259 5952 19323 5956
rect 19339 6012 19403 6016
rect 19339 5956 19343 6012
rect 19343 5956 19399 6012
rect 19399 5956 19403 6012
rect 19339 5952 19403 5956
rect 19419 6012 19483 6016
rect 19419 5956 19423 6012
rect 19423 5956 19479 6012
rect 19479 5956 19483 6012
rect 19419 5952 19483 5956
rect 19499 6012 19563 6016
rect 19499 5956 19503 6012
rect 19503 5956 19559 6012
rect 19559 5956 19563 6012
rect 19499 5952 19563 5956
rect 2757 5468 2821 5472
rect 2757 5412 2761 5468
rect 2761 5412 2817 5468
rect 2817 5412 2821 5468
rect 2757 5408 2821 5412
rect 2837 5468 2901 5472
rect 2837 5412 2841 5468
rect 2841 5412 2897 5468
rect 2897 5412 2901 5468
rect 2837 5408 2901 5412
rect 2917 5468 2981 5472
rect 2917 5412 2921 5468
rect 2921 5412 2977 5468
rect 2977 5412 2981 5468
rect 2917 5408 2981 5412
rect 2997 5468 3061 5472
rect 2997 5412 3001 5468
rect 3001 5412 3057 5468
rect 3057 5412 3061 5468
rect 2997 5408 3061 5412
rect 7472 5468 7536 5472
rect 7472 5412 7476 5468
rect 7476 5412 7532 5468
rect 7532 5412 7536 5468
rect 7472 5408 7536 5412
rect 7552 5468 7616 5472
rect 7552 5412 7556 5468
rect 7556 5412 7612 5468
rect 7612 5412 7616 5468
rect 7552 5408 7616 5412
rect 7632 5468 7696 5472
rect 7632 5412 7636 5468
rect 7636 5412 7692 5468
rect 7692 5412 7696 5468
rect 7632 5408 7696 5412
rect 7712 5468 7776 5472
rect 7712 5412 7716 5468
rect 7716 5412 7772 5468
rect 7772 5412 7776 5468
rect 7712 5408 7776 5412
rect 12187 5468 12251 5472
rect 12187 5412 12191 5468
rect 12191 5412 12247 5468
rect 12247 5412 12251 5468
rect 12187 5408 12251 5412
rect 12267 5468 12331 5472
rect 12267 5412 12271 5468
rect 12271 5412 12327 5468
rect 12327 5412 12331 5468
rect 12267 5408 12331 5412
rect 12347 5468 12411 5472
rect 12347 5412 12351 5468
rect 12351 5412 12407 5468
rect 12407 5412 12411 5468
rect 12347 5408 12411 5412
rect 12427 5468 12491 5472
rect 12427 5412 12431 5468
rect 12431 5412 12487 5468
rect 12487 5412 12491 5468
rect 12427 5408 12491 5412
rect 16902 5468 16966 5472
rect 16902 5412 16906 5468
rect 16906 5412 16962 5468
rect 16962 5412 16966 5468
rect 16902 5408 16966 5412
rect 16982 5468 17046 5472
rect 16982 5412 16986 5468
rect 16986 5412 17042 5468
rect 17042 5412 17046 5468
rect 16982 5408 17046 5412
rect 17062 5468 17126 5472
rect 17062 5412 17066 5468
rect 17066 5412 17122 5468
rect 17122 5412 17126 5468
rect 17062 5408 17126 5412
rect 17142 5468 17206 5472
rect 17142 5412 17146 5468
rect 17146 5412 17202 5468
rect 17202 5412 17206 5468
rect 17142 5408 17206 5412
rect 5114 4924 5178 4928
rect 5114 4868 5118 4924
rect 5118 4868 5174 4924
rect 5174 4868 5178 4924
rect 5114 4864 5178 4868
rect 5194 4924 5258 4928
rect 5194 4868 5198 4924
rect 5198 4868 5254 4924
rect 5254 4868 5258 4924
rect 5194 4864 5258 4868
rect 5274 4924 5338 4928
rect 5274 4868 5278 4924
rect 5278 4868 5334 4924
rect 5334 4868 5338 4924
rect 5274 4864 5338 4868
rect 5354 4924 5418 4928
rect 5354 4868 5358 4924
rect 5358 4868 5414 4924
rect 5414 4868 5418 4924
rect 5354 4864 5418 4868
rect 9829 4924 9893 4928
rect 9829 4868 9833 4924
rect 9833 4868 9889 4924
rect 9889 4868 9893 4924
rect 9829 4864 9893 4868
rect 9909 4924 9973 4928
rect 9909 4868 9913 4924
rect 9913 4868 9969 4924
rect 9969 4868 9973 4924
rect 9909 4864 9973 4868
rect 9989 4924 10053 4928
rect 9989 4868 9993 4924
rect 9993 4868 10049 4924
rect 10049 4868 10053 4924
rect 9989 4864 10053 4868
rect 10069 4924 10133 4928
rect 10069 4868 10073 4924
rect 10073 4868 10129 4924
rect 10129 4868 10133 4924
rect 10069 4864 10133 4868
rect 14544 4924 14608 4928
rect 14544 4868 14548 4924
rect 14548 4868 14604 4924
rect 14604 4868 14608 4924
rect 14544 4864 14608 4868
rect 14624 4924 14688 4928
rect 14624 4868 14628 4924
rect 14628 4868 14684 4924
rect 14684 4868 14688 4924
rect 14624 4864 14688 4868
rect 14704 4924 14768 4928
rect 14704 4868 14708 4924
rect 14708 4868 14764 4924
rect 14764 4868 14768 4924
rect 14704 4864 14768 4868
rect 14784 4924 14848 4928
rect 14784 4868 14788 4924
rect 14788 4868 14844 4924
rect 14844 4868 14848 4924
rect 14784 4864 14848 4868
rect 19259 4924 19323 4928
rect 19259 4868 19263 4924
rect 19263 4868 19319 4924
rect 19319 4868 19323 4924
rect 19259 4864 19323 4868
rect 19339 4924 19403 4928
rect 19339 4868 19343 4924
rect 19343 4868 19399 4924
rect 19399 4868 19403 4924
rect 19339 4864 19403 4868
rect 19419 4924 19483 4928
rect 19419 4868 19423 4924
rect 19423 4868 19479 4924
rect 19479 4868 19483 4924
rect 19419 4864 19483 4868
rect 19499 4924 19563 4928
rect 19499 4868 19503 4924
rect 19503 4868 19559 4924
rect 19559 4868 19563 4924
rect 19499 4864 19563 4868
rect 2757 4380 2821 4384
rect 2757 4324 2761 4380
rect 2761 4324 2817 4380
rect 2817 4324 2821 4380
rect 2757 4320 2821 4324
rect 2837 4380 2901 4384
rect 2837 4324 2841 4380
rect 2841 4324 2897 4380
rect 2897 4324 2901 4380
rect 2837 4320 2901 4324
rect 2917 4380 2981 4384
rect 2917 4324 2921 4380
rect 2921 4324 2977 4380
rect 2977 4324 2981 4380
rect 2917 4320 2981 4324
rect 2997 4380 3061 4384
rect 2997 4324 3001 4380
rect 3001 4324 3057 4380
rect 3057 4324 3061 4380
rect 2997 4320 3061 4324
rect 7472 4380 7536 4384
rect 7472 4324 7476 4380
rect 7476 4324 7532 4380
rect 7532 4324 7536 4380
rect 7472 4320 7536 4324
rect 7552 4380 7616 4384
rect 7552 4324 7556 4380
rect 7556 4324 7612 4380
rect 7612 4324 7616 4380
rect 7552 4320 7616 4324
rect 7632 4380 7696 4384
rect 7632 4324 7636 4380
rect 7636 4324 7692 4380
rect 7692 4324 7696 4380
rect 7632 4320 7696 4324
rect 7712 4380 7776 4384
rect 7712 4324 7716 4380
rect 7716 4324 7772 4380
rect 7772 4324 7776 4380
rect 7712 4320 7776 4324
rect 12187 4380 12251 4384
rect 12187 4324 12191 4380
rect 12191 4324 12247 4380
rect 12247 4324 12251 4380
rect 12187 4320 12251 4324
rect 12267 4380 12331 4384
rect 12267 4324 12271 4380
rect 12271 4324 12327 4380
rect 12327 4324 12331 4380
rect 12267 4320 12331 4324
rect 12347 4380 12411 4384
rect 12347 4324 12351 4380
rect 12351 4324 12407 4380
rect 12407 4324 12411 4380
rect 12347 4320 12411 4324
rect 12427 4380 12491 4384
rect 12427 4324 12431 4380
rect 12431 4324 12487 4380
rect 12487 4324 12491 4380
rect 12427 4320 12491 4324
rect 16902 4380 16966 4384
rect 16902 4324 16906 4380
rect 16906 4324 16962 4380
rect 16962 4324 16966 4380
rect 16902 4320 16966 4324
rect 16982 4380 17046 4384
rect 16982 4324 16986 4380
rect 16986 4324 17042 4380
rect 17042 4324 17046 4380
rect 16982 4320 17046 4324
rect 17062 4380 17126 4384
rect 17062 4324 17066 4380
rect 17066 4324 17122 4380
rect 17122 4324 17126 4380
rect 17062 4320 17126 4324
rect 17142 4380 17206 4384
rect 17142 4324 17146 4380
rect 17146 4324 17202 4380
rect 17202 4324 17206 4380
rect 17142 4320 17206 4324
rect 5114 3836 5178 3840
rect 5114 3780 5118 3836
rect 5118 3780 5174 3836
rect 5174 3780 5178 3836
rect 5114 3776 5178 3780
rect 5194 3836 5258 3840
rect 5194 3780 5198 3836
rect 5198 3780 5254 3836
rect 5254 3780 5258 3836
rect 5194 3776 5258 3780
rect 5274 3836 5338 3840
rect 5274 3780 5278 3836
rect 5278 3780 5334 3836
rect 5334 3780 5338 3836
rect 5274 3776 5338 3780
rect 5354 3836 5418 3840
rect 5354 3780 5358 3836
rect 5358 3780 5414 3836
rect 5414 3780 5418 3836
rect 5354 3776 5418 3780
rect 9829 3836 9893 3840
rect 9829 3780 9833 3836
rect 9833 3780 9889 3836
rect 9889 3780 9893 3836
rect 9829 3776 9893 3780
rect 9909 3836 9973 3840
rect 9909 3780 9913 3836
rect 9913 3780 9969 3836
rect 9969 3780 9973 3836
rect 9909 3776 9973 3780
rect 9989 3836 10053 3840
rect 9989 3780 9993 3836
rect 9993 3780 10049 3836
rect 10049 3780 10053 3836
rect 9989 3776 10053 3780
rect 10069 3836 10133 3840
rect 10069 3780 10073 3836
rect 10073 3780 10129 3836
rect 10129 3780 10133 3836
rect 10069 3776 10133 3780
rect 14544 3836 14608 3840
rect 14544 3780 14548 3836
rect 14548 3780 14604 3836
rect 14604 3780 14608 3836
rect 14544 3776 14608 3780
rect 14624 3836 14688 3840
rect 14624 3780 14628 3836
rect 14628 3780 14684 3836
rect 14684 3780 14688 3836
rect 14624 3776 14688 3780
rect 14704 3836 14768 3840
rect 14704 3780 14708 3836
rect 14708 3780 14764 3836
rect 14764 3780 14768 3836
rect 14704 3776 14768 3780
rect 14784 3836 14848 3840
rect 14784 3780 14788 3836
rect 14788 3780 14844 3836
rect 14844 3780 14848 3836
rect 14784 3776 14848 3780
rect 19259 3836 19323 3840
rect 19259 3780 19263 3836
rect 19263 3780 19319 3836
rect 19319 3780 19323 3836
rect 19259 3776 19323 3780
rect 19339 3836 19403 3840
rect 19339 3780 19343 3836
rect 19343 3780 19399 3836
rect 19399 3780 19403 3836
rect 19339 3776 19403 3780
rect 19419 3836 19483 3840
rect 19419 3780 19423 3836
rect 19423 3780 19479 3836
rect 19479 3780 19483 3836
rect 19419 3776 19483 3780
rect 19499 3836 19563 3840
rect 19499 3780 19503 3836
rect 19503 3780 19559 3836
rect 19559 3780 19563 3836
rect 19499 3776 19563 3780
rect 2757 3292 2821 3296
rect 2757 3236 2761 3292
rect 2761 3236 2817 3292
rect 2817 3236 2821 3292
rect 2757 3232 2821 3236
rect 2837 3292 2901 3296
rect 2837 3236 2841 3292
rect 2841 3236 2897 3292
rect 2897 3236 2901 3292
rect 2837 3232 2901 3236
rect 2917 3292 2981 3296
rect 2917 3236 2921 3292
rect 2921 3236 2977 3292
rect 2977 3236 2981 3292
rect 2917 3232 2981 3236
rect 2997 3292 3061 3296
rect 2997 3236 3001 3292
rect 3001 3236 3057 3292
rect 3057 3236 3061 3292
rect 2997 3232 3061 3236
rect 7472 3292 7536 3296
rect 7472 3236 7476 3292
rect 7476 3236 7532 3292
rect 7532 3236 7536 3292
rect 7472 3232 7536 3236
rect 7552 3292 7616 3296
rect 7552 3236 7556 3292
rect 7556 3236 7612 3292
rect 7612 3236 7616 3292
rect 7552 3232 7616 3236
rect 7632 3292 7696 3296
rect 7632 3236 7636 3292
rect 7636 3236 7692 3292
rect 7692 3236 7696 3292
rect 7632 3232 7696 3236
rect 7712 3292 7776 3296
rect 7712 3236 7716 3292
rect 7716 3236 7772 3292
rect 7772 3236 7776 3292
rect 7712 3232 7776 3236
rect 12187 3292 12251 3296
rect 12187 3236 12191 3292
rect 12191 3236 12247 3292
rect 12247 3236 12251 3292
rect 12187 3232 12251 3236
rect 12267 3292 12331 3296
rect 12267 3236 12271 3292
rect 12271 3236 12327 3292
rect 12327 3236 12331 3292
rect 12267 3232 12331 3236
rect 12347 3292 12411 3296
rect 12347 3236 12351 3292
rect 12351 3236 12407 3292
rect 12407 3236 12411 3292
rect 12347 3232 12411 3236
rect 12427 3292 12491 3296
rect 12427 3236 12431 3292
rect 12431 3236 12487 3292
rect 12487 3236 12491 3292
rect 12427 3232 12491 3236
rect 16902 3292 16966 3296
rect 16902 3236 16906 3292
rect 16906 3236 16962 3292
rect 16962 3236 16966 3292
rect 16902 3232 16966 3236
rect 16982 3292 17046 3296
rect 16982 3236 16986 3292
rect 16986 3236 17042 3292
rect 17042 3236 17046 3292
rect 16982 3232 17046 3236
rect 17062 3292 17126 3296
rect 17062 3236 17066 3292
rect 17066 3236 17122 3292
rect 17122 3236 17126 3292
rect 17062 3232 17126 3236
rect 17142 3292 17206 3296
rect 17142 3236 17146 3292
rect 17146 3236 17202 3292
rect 17202 3236 17206 3292
rect 17142 3232 17206 3236
rect 5114 2748 5178 2752
rect 5114 2692 5118 2748
rect 5118 2692 5174 2748
rect 5174 2692 5178 2748
rect 5114 2688 5178 2692
rect 5194 2748 5258 2752
rect 5194 2692 5198 2748
rect 5198 2692 5254 2748
rect 5254 2692 5258 2748
rect 5194 2688 5258 2692
rect 5274 2748 5338 2752
rect 5274 2692 5278 2748
rect 5278 2692 5334 2748
rect 5334 2692 5338 2748
rect 5274 2688 5338 2692
rect 5354 2748 5418 2752
rect 5354 2692 5358 2748
rect 5358 2692 5414 2748
rect 5414 2692 5418 2748
rect 5354 2688 5418 2692
rect 9829 2748 9893 2752
rect 9829 2692 9833 2748
rect 9833 2692 9889 2748
rect 9889 2692 9893 2748
rect 9829 2688 9893 2692
rect 9909 2748 9973 2752
rect 9909 2692 9913 2748
rect 9913 2692 9969 2748
rect 9969 2692 9973 2748
rect 9909 2688 9973 2692
rect 9989 2748 10053 2752
rect 9989 2692 9993 2748
rect 9993 2692 10049 2748
rect 10049 2692 10053 2748
rect 9989 2688 10053 2692
rect 10069 2748 10133 2752
rect 10069 2692 10073 2748
rect 10073 2692 10129 2748
rect 10129 2692 10133 2748
rect 10069 2688 10133 2692
rect 14544 2748 14608 2752
rect 14544 2692 14548 2748
rect 14548 2692 14604 2748
rect 14604 2692 14608 2748
rect 14544 2688 14608 2692
rect 14624 2748 14688 2752
rect 14624 2692 14628 2748
rect 14628 2692 14684 2748
rect 14684 2692 14688 2748
rect 14624 2688 14688 2692
rect 14704 2748 14768 2752
rect 14704 2692 14708 2748
rect 14708 2692 14764 2748
rect 14764 2692 14768 2748
rect 14704 2688 14768 2692
rect 14784 2748 14848 2752
rect 14784 2692 14788 2748
rect 14788 2692 14844 2748
rect 14844 2692 14848 2748
rect 14784 2688 14848 2692
rect 19259 2748 19323 2752
rect 19259 2692 19263 2748
rect 19263 2692 19319 2748
rect 19319 2692 19323 2748
rect 19259 2688 19323 2692
rect 19339 2748 19403 2752
rect 19339 2692 19343 2748
rect 19343 2692 19399 2748
rect 19399 2692 19403 2748
rect 19339 2688 19403 2692
rect 19419 2748 19483 2752
rect 19419 2692 19423 2748
rect 19423 2692 19479 2748
rect 19479 2692 19483 2748
rect 19419 2688 19483 2692
rect 19499 2748 19563 2752
rect 19499 2692 19503 2748
rect 19503 2692 19559 2748
rect 19559 2692 19563 2748
rect 19499 2688 19563 2692
rect 2757 2204 2821 2208
rect 2757 2148 2761 2204
rect 2761 2148 2817 2204
rect 2817 2148 2821 2204
rect 2757 2144 2821 2148
rect 2837 2204 2901 2208
rect 2837 2148 2841 2204
rect 2841 2148 2897 2204
rect 2897 2148 2901 2204
rect 2837 2144 2901 2148
rect 2917 2204 2981 2208
rect 2917 2148 2921 2204
rect 2921 2148 2977 2204
rect 2977 2148 2981 2204
rect 2917 2144 2981 2148
rect 2997 2204 3061 2208
rect 2997 2148 3001 2204
rect 3001 2148 3057 2204
rect 3057 2148 3061 2204
rect 2997 2144 3061 2148
rect 7472 2204 7536 2208
rect 7472 2148 7476 2204
rect 7476 2148 7532 2204
rect 7532 2148 7536 2204
rect 7472 2144 7536 2148
rect 7552 2204 7616 2208
rect 7552 2148 7556 2204
rect 7556 2148 7612 2204
rect 7612 2148 7616 2204
rect 7552 2144 7616 2148
rect 7632 2204 7696 2208
rect 7632 2148 7636 2204
rect 7636 2148 7692 2204
rect 7692 2148 7696 2204
rect 7632 2144 7696 2148
rect 7712 2204 7776 2208
rect 7712 2148 7716 2204
rect 7716 2148 7772 2204
rect 7772 2148 7776 2204
rect 7712 2144 7776 2148
rect 12187 2204 12251 2208
rect 12187 2148 12191 2204
rect 12191 2148 12247 2204
rect 12247 2148 12251 2204
rect 12187 2144 12251 2148
rect 12267 2204 12331 2208
rect 12267 2148 12271 2204
rect 12271 2148 12327 2204
rect 12327 2148 12331 2204
rect 12267 2144 12331 2148
rect 12347 2204 12411 2208
rect 12347 2148 12351 2204
rect 12351 2148 12407 2204
rect 12407 2148 12411 2204
rect 12347 2144 12411 2148
rect 12427 2204 12491 2208
rect 12427 2148 12431 2204
rect 12431 2148 12487 2204
rect 12487 2148 12491 2204
rect 12427 2144 12491 2148
rect 16902 2204 16966 2208
rect 16902 2148 16906 2204
rect 16906 2148 16962 2204
rect 16962 2148 16966 2204
rect 16902 2144 16966 2148
rect 16982 2204 17046 2208
rect 16982 2148 16986 2204
rect 16986 2148 17042 2204
rect 17042 2148 17046 2204
rect 16982 2144 17046 2148
rect 17062 2204 17126 2208
rect 17062 2148 17066 2204
rect 17066 2148 17122 2204
rect 17122 2148 17126 2204
rect 17062 2144 17126 2148
rect 17142 2204 17206 2208
rect 17142 2148 17146 2204
rect 17146 2148 17202 2204
rect 17202 2148 17206 2204
rect 17142 2144 17206 2148
rect 5114 1660 5178 1664
rect 5114 1604 5118 1660
rect 5118 1604 5174 1660
rect 5174 1604 5178 1660
rect 5114 1600 5178 1604
rect 5194 1660 5258 1664
rect 5194 1604 5198 1660
rect 5198 1604 5254 1660
rect 5254 1604 5258 1660
rect 5194 1600 5258 1604
rect 5274 1660 5338 1664
rect 5274 1604 5278 1660
rect 5278 1604 5334 1660
rect 5334 1604 5338 1660
rect 5274 1600 5338 1604
rect 5354 1660 5418 1664
rect 5354 1604 5358 1660
rect 5358 1604 5414 1660
rect 5414 1604 5418 1660
rect 5354 1600 5418 1604
rect 9829 1660 9893 1664
rect 9829 1604 9833 1660
rect 9833 1604 9889 1660
rect 9889 1604 9893 1660
rect 9829 1600 9893 1604
rect 9909 1660 9973 1664
rect 9909 1604 9913 1660
rect 9913 1604 9969 1660
rect 9969 1604 9973 1660
rect 9909 1600 9973 1604
rect 9989 1660 10053 1664
rect 9989 1604 9993 1660
rect 9993 1604 10049 1660
rect 10049 1604 10053 1660
rect 9989 1600 10053 1604
rect 10069 1660 10133 1664
rect 10069 1604 10073 1660
rect 10073 1604 10129 1660
rect 10129 1604 10133 1660
rect 10069 1600 10133 1604
rect 14544 1660 14608 1664
rect 14544 1604 14548 1660
rect 14548 1604 14604 1660
rect 14604 1604 14608 1660
rect 14544 1600 14608 1604
rect 14624 1660 14688 1664
rect 14624 1604 14628 1660
rect 14628 1604 14684 1660
rect 14684 1604 14688 1660
rect 14624 1600 14688 1604
rect 14704 1660 14768 1664
rect 14704 1604 14708 1660
rect 14708 1604 14764 1660
rect 14764 1604 14768 1660
rect 14704 1600 14768 1604
rect 14784 1660 14848 1664
rect 14784 1604 14788 1660
rect 14788 1604 14844 1660
rect 14844 1604 14848 1660
rect 14784 1600 14848 1604
rect 19259 1660 19323 1664
rect 19259 1604 19263 1660
rect 19263 1604 19319 1660
rect 19319 1604 19323 1660
rect 19259 1600 19323 1604
rect 19339 1660 19403 1664
rect 19339 1604 19343 1660
rect 19343 1604 19399 1660
rect 19399 1604 19403 1660
rect 19339 1600 19403 1604
rect 19419 1660 19483 1664
rect 19419 1604 19423 1660
rect 19423 1604 19479 1660
rect 19479 1604 19483 1660
rect 19419 1600 19483 1604
rect 19499 1660 19563 1664
rect 19499 1604 19503 1660
rect 19503 1604 19559 1660
rect 19559 1604 19563 1660
rect 19499 1600 19563 1604
rect 2757 1116 2821 1120
rect 2757 1060 2761 1116
rect 2761 1060 2817 1116
rect 2817 1060 2821 1116
rect 2757 1056 2821 1060
rect 2837 1116 2901 1120
rect 2837 1060 2841 1116
rect 2841 1060 2897 1116
rect 2897 1060 2901 1116
rect 2837 1056 2901 1060
rect 2917 1116 2981 1120
rect 2917 1060 2921 1116
rect 2921 1060 2977 1116
rect 2977 1060 2981 1116
rect 2917 1056 2981 1060
rect 2997 1116 3061 1120
rect 2997 1060 3001 1116
rect 3001 1060 3057 1116
rect 3057 1060 3061 1116
rect 2997 1056 3061 1060
rect 7472 1116 7536 1120
rect 7472 1060 7476 1116
rect 7476 1060 7532 1116
rect 7532 1060 7536 1116
rect 7472 1056 7536 1060
rect 7552 1116 7616 1120
rect 7552 1060 7556 1116
rect 7556 1060 7612 1116
rect 7612 1060 7616 1116
rect 7552 1056 7616 1060
rect 7632 1116 7696 1120
rect 7632 1060 7636 1116
rect 7636 1060 7692 1116
rect 7692 1060 7696 1116
rect 7632 1056 7696 1060
rect 7712 1116 7776 1120
rect 7712 1060 7716 1116
rect 7716 1060 7772 1116
rect 7772 1060 7776 1116
rect 7712 1056 7776 1060
rect 12187 1116 12251 1120
rect 12187 1060 12191 1116
rect 12191 1060 12247 1116
rect 12247 1060 12251 1116
rect 12187 1056 12251 1060
rect 12267 1116 12331 1120
rect 12267 1060 12271 1116
rect 12271 1060 12327 1116
rect 12327 1060 12331 1116
rect 12267 1056 12331 1060
rect 12347 1116 12411 1120
rect 12347 1060 12351 1116
rect 12351 1060 12407 1116
rect 12407 1060 12411 1116
rect 12347 1056 12411 1060
rect 12427 1116 12491 1120
rect 12427 1060 12431 1116
rect 12431 1060 12487 1116
rect 12487 1060 12491 1116
rect 12427 1056 12491 1060
rect 16902 1116 16966 1120
rect 16902 1060 16906 1116
rect 16906 1060 16962 1116
rect 16962 1060 16966 1116
rect 16902 1056 16966 1060
rect 16982 1116 17046 1120
rect 16982 1060 16986 1116
rect 16986 1060 17042 1116
rect 17042 1060 17046 1116
rect 16982 1056 17046 1060
rect 17062 1116 17126 1120
rect 17062 1060 17066 1116
rect 17066 1060 17122 1116
rect 17122 1060 17126 1116
rect 17062 1056 17126 1060
rect 17142 1116 17206 1120
rect 17142 1060 17146 1116
rect 17146 1060 17202 1116
rect 17202 1060 17206 1116
rect 17142 1056 17206 1060
rect 5114 572 5178 576
rect 5114 516 5118 572
rect 5118 516 5174 572
rect 5174 516 5178 572
rect 5114 512 5178 516
rect 5194 572 5258 576
rect 5194 516 5198 572
rect 5198 516 5254 572
rect 5254 516 5258 572
rect 5194 512 5258 516
rect 5274 572 5338 576
rect 5274 516 5278 572
rect 5278 516 5334 572
rect 5334 516 5338 572
rect 5274 512 5338 516
rect 5354 572 5418 576
rect 5354 516 5358 572
rect 5358 516 5414 572
rect 5414 516 5418 572
rect 5354 512 5418 516
rect 9829 572 9893 576
rect 9829 516 9833 572
rect 9833 516 9889 572
rect 9889 516 9893 572
rect 9829 512 9893 516
rect 9909 572 9973 576
rect 9909 516 9913 572
rect 9913 516 9969 572
rect 9969 516 9973 572
rect 9909 512 9973 516
rect 9989 572 10053 576
rect 9989 516 9993 572
rect 9993 516 10049 572
rect 10049 516 10053 572
rect 9989 512 10053 516
rect 10069 572 10133 576
rect 10069 516 10073 572
rect 10073 516 10129 572
rect 10129 516 10133 572
rect 10069 512 10133 516
rect 14544 572 14608 576
rect 14544 516 14548 572
rect 14548 516 14604 572
rect 14604 516 14608 572
rect 14544 512 14608 516
rect 14624 572 14688 576
rect 14624 516 14628 572
rect 14628 516 14684 572
rect 14684 516 14688 572
rect 14624 512 14688 516
rect 14704 572 14768 576
rect 14704 516 14708 572
rect 14708 516 14764 572
rect 14764 516 14768 572
rect 14704 512 14768 516
rect 14784 572 14848 576
rect 14784 516 14788 572
rect 14788 516 14844 572
rect 14844 516 14848 572
rect 14784 512 14848 516
rect 19259 572 19323 576
rect 19259 516 19263 572
rect 19263 516 19319 572
rect 19319 516 19323 572
rect 19259 512 19323 516
rect 19339 572 19403 576
rect 19339 516 19343 572
rect 19343 516 19399 572
rect 19399 516 19403 572
rect 19339 512 19403 516
rect 19419 572 19483 576
rect 19419 516 19423 572
rect 19423 516 19479 572
rect 19479 516 19483 572
rect 19419 512 19483 516
rect 19499 572 19563 576
rect 19499 516 19503 572
rect 19503 516 19559 572
rect 19559 516 19563 572
rect 19499 512 19563 516
<< metal4 >>
rect 2749 18528 3069 19088
rect 2749 18464 2757 18528
rect 2821 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3069 18528
rect 2749 17440 3069 18464
rect 2749 17376 2757 17440
rect 2821 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3069 17440
rect 2749 16352 3069 17376
rect 2749 16288 2757 16352
rect 2821 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3069 16352
rect 2749 15264 3069 16288
rect 2749 15200 2757 15264
rect 2821 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3069 15264
rect 2749 14176 3069 15200
rect 2749 14112 2757 14176
rect 2821 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3069 14176
rect 2749 13088 3069 14112
rect 2749 13024 2757 13088
rect 2821 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3069 13088
rect 2749 12000 3069 13024
rect 2749 11936 2757 12000
rect 2821 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3069 12000
rect 2749 10912 3069 11936
rect 2749 10848 2757 10912
rect 2821 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3069 10912
rect 2749 9824 3069 10848
rect 2749 9760 2757 9824
rect 2821 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3069 9824
rect 2749 8736 3069 9760
rect 2749 8672 2757 8736
rect 2821 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3069 8736
rect 2749 7648 3069 8672
rect 2749 7584 2757 7648
rect 2821 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3069 7648
rect 2749 6560 3069 7584
rect 2749 6496 2757 6560
rect 2821 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3069 6560
rect 2749 5472 3069 6496
rect 2749 5408 2757 5472
rect 2821 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3069 5472
rect 2749 4384 3069 5408
rect 2749 4320 2757 4384
rect 2821 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3069 4384
rect 2749 3296 3069 4320
rect 2749 3232 2757 3296
rect 2821 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3069 3296
rect 2749 2208 3069 3232
rect 2749 2144 2757 2208
rect 2821 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3069 2208
rect 2749 1120 3069 2144
rect 2749 1056 2757 1120
rect 2821 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3069 1120
rect 2749 496 3069 1056
rect 5106 19072 5426 19088
rect 5106 19008 5114 19072
rect 5178 19008 5194 19072
rect 5258 19008 5274 19072
rect 5338 19008 5354 19072
rect 5418 19008 5426 19072
rect 5106 17984 5426 19008
rect 5106 17920 5114 17984
rect 5178 17920 5194 17984
rect 5258 17920 5274 17984
rect 5338 17920 5354 17984
rect 5418 17920 5426 17984
rect 5106 16896 5426 17920
rect 5106 16832 5114 16896
rect 5178 16832 5194 16896
rect 5258 16832 5274 16896
rect 5338 16832 5354 16896
rect 5418 16832 5426 16896
rect 5106 15808 5426 16832
rect 5106 15744 5114 15808
rect 5178 15744 5194 15808
rect 5258 15744 5274 15808
rect 5338 15744 5354 15808
rect 5418 15744 5426 15808
rect 5106 14720 5426 15744
rect 5106 14656 5114 14720
rect 5178 14656 5194 14720
rect 5258 14656 5274 14720
rect 5338 14656 5354 14720
rect 5418 14656 5426 14720
rect 5106 13632 5426 14656
rect 5106 13568 5114 13632
rect 5178 13568 5194 13632
rect 5258 13568 5274 13632
rect 5338 13568 5354 13632
rect 5418 13568 5426 13632
rect 5106 12544 5426 13568
rect 5106 12480 5114 12544
rect 5178 12480 5194 12544
rect 5258 12480 5274 12544
rect 5338 12480 5354 12544
rect 5418 12480 5426 12544
rect 5106 11456 5426 12480
rect 5106 11392 5114 11456
rect 5178 11392 5194 11456
rect 5258 11392 5274 11456
rect 5338 11392 5354 11456
rect 5418 11392 5426 11456
rect 5106 10368 5426 11392
rect 5106 10304 5114 10368
rect 5178 10304 5194 10368
rect 5258 10304 5274 10368
rect 5338 10304 5354 10368
rect 5418 10304 5426 10368
rect 5106 9280 5426 10304
rect 5106 9216 5114 9280
rect 5178 9216 5194 9280
rect 5258 9216 5274 9280
rect 5338 9216 5354 9280
rect 5418 9216 5426 9280
rect 5106 8192 5426 9216
rect 5106 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5354 8192
rect 5418 8128 5426 8192
rect 5106 7104 5426 8128
rect 5106 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5354 7104
rect 5418 7040 5426 7104
rect 5106 6016 5426 7040
rect 5106 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5354 6016
rect 5418 5952 5426 6016
rect 5106 4928 5426 5952
rect 5106 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5354 4928
rect 5418 4864 5426 4928
rect 5106 3840 5426 4864
rect 5106 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5354 3840
rect 5418 3776 5426 3840
rect 5106 2752 5426 3776
rect 5106 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5354 2752
rect 5418 2688 5426 2752
rect 5106 1664 5426 2688
rect 5106 1600 5114 1664
rect 5178 1600 5194 1664
rect 5258 1600 5274 1664
rect 5338 1600 5354 1664
rect 5418 1600 5426 1664
rect 5106 576 5426 1600
rect 5106 512 5114 576
rect 5178 512 5194 576
rect 5258 512 5274 576
rect 5338 512 5354 576
rect 5418 512 5426 576
rect 5106 496 5426 512
rect 7464 18528 7784 19088
rect 7464 18464 7472 18528
rect 7536 18464 7552 18528
rect 7616 18464 7632 18528
rect 7696 18464 7712 18528
rect 7776 18464 7784 18528
rect 7464 17440 7784 18464
rect 7464 17376 7472 17440
rect 7536 17376 7552 17440
rect 7616 17376 7632 17440
rect 7696 17376 7712 17440
rect 7776 17376 7784 17440
rect 7464 16352 7784 17376
rect 7464 16288 7472 16352
rect 7536 16288 7552 16352
rect 7616 16288 7632 16352
rect 7696 16288 7712 16352
rect 7776 16288 7784 16352
rect 7464 15264 7784 16288
rect 7464 15200 7472 15264
rect 7536 15200 7552 15264
rect 7616 15200 7632 15264
rect 7696 15200 7712 15264
rect 7776 15200 7784 15264
rect 7464 14176 7784 15200
rect 7464 14112 7472 14176
rect 7536 14112 7552 14176
rect 7616 14112 7632 14176
rect 7696 14112 7712 14176
rect 7776 14112 7784 14176
rect 7464 13088 7784 14112
rect 7464 13024 7472 13088
rect 7536 13024 7552 13088
rect 7616 13024 7632 13088
rect 7696 13024 7712 13088
rect 7776 13024 7784 13088
rect 7464 12000 7784 13024
rect 7464 11936 7472 12000
rect 7536 11936 7552 12000
rect 7616 11936 7632 12000
rect 7696 11936 7712 12000
rect 7776 11936 7784 12000
rect 7464 10912 7784 11936
rect 7464 10848 7472 10912
rect 7536 10848 7552 10912
rect 7616 10848 7632 10912
rect 7696 10848 7712 10912
rect 7776 10848 7784 10912
rect 7464 9824 7784 10848
rect 7464 9760 7472 9824
rect 7536 9760 7552 9824
rect 7616 9760 7632 9824
rect 7696 9760 7712 9824
rect 7776 9760 7784 9824
rect 7464 8736 7784 9760
rect 7464 8672 7472 8736
rect 7536 8672 7552 8736
rect 7616 8672 7632 8736
rect 7696 8672 7712 8736
rect 7776 8672 7784 8736
rect 7464 7648 7784 8672
rect 7464 7584 7472 7648
rect 7536 7584 7552 7648
rect 7616 7584 7632 7648
rect 7696 7584 7712 7648
rect 7776 7584 7784 7648
rect 7464 6560 7784 7584
rect 7464 6496 7472 6560
rect 7536 6496 7552 6560
rect 7616 6496 7632 6560
rect 7696 6496 7712 6560
rect 7776 6496 7784 6560
rect 7464 5472 7784 6496
rect 7464 5408 7472 5472
rect 7536 5408 7552 5472
rect 7616 5408 7632 5472
rect 7696 5408 7712 5472
rect 7776 5408 7784 5472
rect 7464 4384 7784 5408
rect 7464 4320 7472 4384
rect 7536 4320 7552 4384
rect 7616 4320 7632 4384
rect 7696 4320 7712 4384
rect 7776 4320 7784 4384
rect 7464 3296 7784 4320
rect 7464 3232 7472 3296
rect 7536 3232 7552 3296
rect 7616 3232 7632 3296
rect 7696 3232 7712 3296
rect 7776 3232 7784 3296
rect 7464 2208 7784 3232
rect 7464 2144 7472 2208
rect 7536 2144 7552 2208
rect 7616 2144 7632 2208
rect 7696 2144 7712 2208
rect 7776 2144 7784 2208
rect 7464 1120 7784 2144
rect 7464 1056 7472 1120
rect 7536 1056 7552 1120
rect 7616 1056 7632 1120
rect 7696 1056 7712 1120
rect 7776 1056 7784 1120
rect 7464 496 7784 1056
rect 9821 19072 10141 19088
rect 9821 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10069 19072
rect 10133 19008 10141 19072
rect 9821 17984 10141 19008
rect 9821 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10069 17984
rect 10133 17920 10141 17984
rect 9821 16896 10141 17920
rect 9821 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10069 16896
rect 10133 16832 10141 16896
rect 9821 15808 10141 16832
rect 9821 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10069 15808
rect 10133 15744 10141 15808
rect 9821 14720 10141 15744
rect 9821 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10069 14720
rect 10133 14656 10141 14720
rect 9821 13632 10141 14656
rect 9821 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10069 13632
rect 10133 13568 10141 13632
rect 9821 12544 10141 13568
rect 9821 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10069 12544
rect 10133 12480 10141 12544
rect 9821 11456 10141 12480
rect 9821 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10069 11456
rect 10133 11392 10141 11456
rect 9821 10368 10141 11392
rect 9821 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10069 10368
rect 10133 10304 10141 10368
rect 9821 9280 10141 10304
rect 9821 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10069 9280
rect 10133 9216 10141 9280
rect 9821 8192 10141 9216
rect 9821 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10069 8192
rect 10133 8128 10141 8192
rect 9821 7104 10141 8128
rect 9821 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10069 7104
rect 10133 7040 10141 7104
rect 9821 6016 10141 7040
rect 9821 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10069 6016
rect 10133 5952 10141 6016
rect 9821 4928 10141 5952
rect 9821 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10069 4928
rect 10133 4864 10141 4928
rect 9821 3840 10141 4864
rect 9821 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10069 3840
rect 10133 3776 10141 3840
rect 9821 2752 10141 3776
rect 9821 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10069 2752
rect 10133 2688 10141 2752
rect 9821 1664 10141 2688
rect 9821 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10069 1664
rect 10133 1600 10141 1664
rect 9821 576 10141 1600
rect 9821 512 9829 576
rect 9893 512 9909 576
rect 9973 512 9989 576
rect 10053 512 10069 576
rect 10133 512 10141 576
rect 9821 496 10141 512
rect 12179 18528 12499 19088
rect 12179 18464 12187 18528
rect 12251 18464 12267 18528
rect 12331 18464 12347 18528
rect 12411 18464 12427 18528
rect 12491 18464 12499 18528
rect 12179 17440 12499 18464
rect 12179 17376 12187 17440
rect 12251 17376 12267 17440
rect 12331 17376 12347 17440
rect 12411 17376 12427 17440
rect 12491 17376 12499 17440
rect 12179 16352 12499 17376
rect 12179 16288 12187 16352
rect 12251 16288 12267 16352
rect 12331 16288 12347 16352
rect 12411 16288 12427 16352
rect 12491 16288 12499 16352
rect 12179 15264 12499 16288
rect 12179 15200 12187 15264
rect 12251 15200 12267 15264
rect 12331 15200 12347 15264
rect 12411 15200 12427 15264
rect 12491 15200 12499 15264
rect 12179 14176 12499 15200
rect 12179 14112 12187 14176
rect 12251 14112 12267 14176
rect 12331 14112 12347 14176
rect 12411 14112 12427 14176
rect 12491 14112 12499 14176
rect 12179 13088 12499 14112
rect 12179 13024 12187 13088
rect 12251 13024 12267 13088
rect 12331 13024 12347 13088
rect 12411 13024 12427 13088
rect 12491 13024 12499 13088
rect 12179 12000 12499 13024
rect 12179 11936 12187 12000
rect 12251 11936 12267 12000
rect 12331 11936 12347 12000
rect 12411 11936 12427 12000
rect 12491 11936 12499 12000
rect 12179 10912 12499 11936
rect 12179 10848 12187 10912
rect 12251 10848 12267 10912
rect 12331 10848 12347 10912
rect 12411 10848 12427 10912
rect 12491 10848 12499 10912
rect 12179 9824 12499 10848
rect 12179 9760 12187 9824
rect 12251 9760 12267 9824
rect 12331 9760 12347 9824
rect 12411 9760 12427 9824
rect 12491 9760 12499 9824
rect 12179 8736 12499 9760
rect 12179 8672 12187 8736
rect 12251 8672 12267 8736
rect 12331 8672 12347 8736
rect 12411 8672 12427 8736
rect 12491 8672 12499 8736
rect 12179 7648 12499 8672
rect 12179 7584 12187 7648
rect 12251 7584 12267 7648
rect 12331 7584 12347 7648
rect 12411 7584 12427 7648
rect 12491 7584 12499 7648
rect 12179 6560 12499 7584
rect 12179 6496 12187 6560
rect 12251 6496 12267 6560
rect 12331 6496 12347 6560
rect 12411 6496 12427 6560
rect 12491 6496 12499 6560
rect 12179 5472 12499 6496
rect 12179 5408 12187 5472
rect 12251 5408 12267 5472
rect 12331 5408 12347 5472
rect 12411 5408 12427 5472
rect 12491 5408 12499 5472
rect 12179 4384 12499 5408
rect 12179 4320 12187 4384
rect 12251 4320 12267 4384
rect 12331 4320 12347 4384
rect 12411 4320 12427 4384
rect 12491 4320 12499 4384
rect 12179 3296 12499 4320
rect 12179 3232 12187 3296
rect 12251 3232 12267 3296
rect 12331 3232 12347 3296
rect 12411 3232 12427 3296
rect 12491 3232 12499 3296
rect 12179 2208 12499 3232
rect 12179 2144 12187 2208
rect 12251 2144 12267 2208
rect 12331 2144 12347 2208
rect 12411 2144 12427 2208
rect 12491 2144 12499 2208
rect 12179 1120 12499 2144
rect 12179 1056 12187 1120
rect 12251 1056 12267 1120
rect 12331 1056 12347 1120
rect 12411 1056 12427 1120
rect 12491 1056 12499 1120
rect 12179 496 12499 1056
rect 14536 19072 14856 19088
rect 14536 19008 14544 19072
rect 14608 19008 14624 19072
rect 14688 19008 14704 19072
rect 14768 19008 14784 19072
rect 14848 19008 14856 19072
rect 14536 17984 14856 19008
rect 14536 17920 14544 17984
rect 14608 17920 14624 17984
rect 14688 17920 14704 17984
rect 14768 17920 14784 17984
rect 14848 17920 14856 17984
rect 14536 16896 14856 17920
rect 14536 16832 14544 16896
rect 14608 16832 14624 16896
rect 14688 16832 14704 16896
rect 14768 16832 14784 16896
rect 14848 16832 14856 16896
rect 14536 15808 14856 16832
rect 14536 15744 14544 15808
rect 14608 15744 14624 15808
rect 14688 15744 14704 15808
rect 14768 15744 14784 15808
rect 14848 15744 14856 15808
rect 14536 14720 14856 15744
rect 14536 14656 14544 14720
rect 14608 14656 14624 14720
rect 14688 14656 14704 14720
rect 14768 14656 14784 14720
rect 14848 14656 14856 14720
rect 14536 13632 14856 14656
rect 14536 13568 14544 13632
rect 14608 13568 14624 13632
rect 14688 13568 14704 13632
rect 14768 13568 14784 13632
rect 14848 13568 14856 13632
rect 14536 12544 14856 13568
rect 14536 12480 14544 12544
rect 14608 12480 14624 12544
rect 14688 12480 14704 12544
rect 14768 12480 14784 12544
rect 14848 12480 14856 12544
rect 14536 11456 14856 12480
rect 14536 11392 14544 11456
rect 14608 11392 14624 11456
rect 14688 11392 14704 11456
rect 14768 11392 14784 11456
rect 14848 11392 14856 11456
rect 14536 10368 14856 11392
rect 14536 10304 14544 10368
rect 14608 10304 14624 10368
rect 14688 10304 14704 10368
rect 14768 10304 14784 10368
rect 14848 10304 14856 10368
rect 14536 9280 14856 10304
rect 14536 9216 14544 9280
rect 14608 9216 14624 9280
rect 14688 9216 14704 9280
rect 14768 9216 14784 9280
rect 14848 9216 14856 9280
rect 14536 8192 14856 9216
rect 14536 8128 14544 8192
rect 14608 8128 14624 8192
rect 14688 8128 14704 8192
rect 14768 8128 14784 8192
rect 14848 8128 14856 8192
rect 14536 7104 14856 8128
rect 14536 7040 14544 7104
rect 14608 7040 14624 7104
rect 14688 7040 14704 7104
rect 14768 7040 14784 7104
rect 14848 7040 14856 7104
rect 14536 6016 14856 7040
rect 14536 5952 14544 6016
rect 14608 5952 14624 6016
rect 14688 5952 14704 6016
rect 14768 5952 14784 6016
rect 14848 5952 14856 6016
rect 14536 4928 14856 5952
rect 14536 4864 14544 4928
rect 14608 4864 14624 4928
rect 14688 4864 14704 4928
rect 14768 4864 14784 4928
rect 14848 4864 14856 4928
rect 14536 3840 14856 4864
rect 14536 3776 14544 3840
rect 14608 3776 14624 3840
rect 14688 3776 14704 3840
rect 14768 3776 14784 3840
rect 14848 3776 14856 3840
rect 14536 2752 14856 3776
rect 14536 2688 14544 2752
rect 14608 2688 14624 2752
rect 14688 2688 14704 2752
rect 14768 2688 14784 2752
rect 14848 2688 14856 2752
rect 14536 1664 14856 2688
rect 14536 1600 14544 1664
rect 14608 1600 14624 1664
rect 14688 1600 14704 1664
rect 14768 1600 14784 1664
rect 14848 1600 14856 1664
rect 14536 576 14856 1600
rect 14536 512 14544 576
rect 14608 512 14624 576
rect 14688 512 14704 576
rect 14768 512 14784 576
rect 14848 512 14856 576
rect 14536 496 14856 512
rect 16894 18528 17214 19088
rect 16894 18464 16902 18528
rect 16966 18464 16982 18528
rect 17046 18464 17062 18528
rect 17126 18464 17142 18528
rect 17206 18464 17214 18528
rect 16894 17440 17214 18464
rect 16894 17376 16902 17440
rect 16966 17376 16982 17440
rect 17046 17376 17062 17440
rect 17126 17376 17142 17440
rect 17206 17376 17214 17440
rect 16894 16352 17214 17376
rect 16894 16288 16902 16352
rect 16966 16288 16982 16352
rect 17046 16288 17062 16352
rect 17126 16288 17142 16352
rect 17206 16288 17214 16352
rect 16894 15264 17214 16288
rect 16894 15200 16902 15264
rect 16966 15200 16982 15264
rect 17046 15200 17062 15264
rect 17126 15200 17142 15264
rect 17206 15200 17214 15264
rect 16894 14176 17214 15200
rect 16894 14112 16902 14176
rect 16966 14112 16982 14176
rect 17046 14112 17062 14176
rect 17126 14112 17142 14176
rect 17206 14112 17214 14176
rect 16894 13088 17214 14112
rect 16894 13024 16902 13088
rect 16966 13024 16982 13088
rect 17046 13024 17062 13088
rect 17126 13024 17142 13088
rect 17206 13024 17214 13088
rect 16894 12000 17214 13024
rect 16894 11936 16902 12000
rect 16966 11936 16982 12000
rect 17046 11936 17062 12000
rect 17126 11936 17142 12000
rect 17206 11936 17214 12000
rect 16894 10912 17214 11936
rect 16894 10848 16902 10912
rect 16966 10848 16982 10912
rect 17046 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17214 10912
rect 16894 9824 17214 10848
rect 16894 9760 16902 9824
rect 16966 9760 16982 9824
rect 17046 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17214 9824
rect 16894 8736 17214 9760
rect 16894 8672 16902 8736
rect 16966 8672 16982 8736
rect 17046 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17214 8736
rect 16894 7648 17214 8672
rect 16894 7584 16902 7648
rect 16966 7584 16982 7648
rect 17046 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17214 7648
rect 16894 6560 17214 7584
rect 16894 6496 16902 6560
rect 16966 6496 16982 6560
rect 17046 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17214 6560
rect 16894 5472 17214 6496
rect 16894 5408 16902 5472
rect 16966 5408 16982 5472
rect 17046 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17214 5472
rect 16894 4384 17214 5408
rect 16894 4320 16902 4384
rect 16966 4320 16982 4384
rect 17046 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17214 4384
rect 16894 3296 17214 4320
rect 16894 3232 16902 3296
rect 16966 3232 16982 3296
rect 17046 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17214 3296
rect 16894 2208 17214 3232
rect 16894 2144 16902 2208
rect 16966 2144 16982 2208
rect 17046 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17214 2208
rect 16894 1120 17214 2144
rect 16894 1056 16902 1120
rect 16966 1056 16982 1120
rect 17046 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17214 1120
rect 16894 496 17214 1056
rect 19251 19072 19571 19088
rect 19251 19008 19259 19072
rect 19323 19008 19339 19072
rect 19403 19008 19419 19072
rect 19483 19008 19499 19072
rect 19563 19008 19571 19072
rect 19251 17984 19571 19008
rect 19251 17920 19259 17984
rect 19323 17920 19339 17984
rect 19403 17920 19419 17984
rect 19483 17920 19499 17984
rect 19563 17920 19571 17984
rect 19251 16896 19571 17920
rect 19251 16832 19259 16896
rect 19323 16832 19339 16896
rect 19403 16832 19419 16896
rect 19483 16832 19499 16896
rect 19563 16832 19571 16896
rect 19251 15808 19571 16832
rect 19251 15744 19259 15808
rect 19323 15744 19339 15808
rect 19403 15744 19419 15808
rect 19483 15744 19499 15808
rect 19563 15744 19571 15808
rect 19251 14720 19571 15744
rect 19251 14656 19259 14720
rect 19323 14656 19339 14720
rect 19403 14656 19419 14720
rect 19483 14656 19499 14720
rect 19563 14656 19571 14720
rect 19251 13632 19571 14656
rect 19251 13568 19259 13632
rect 19323 13568 19339 13632
rect 19403 13568 19419 13632
rect 19483 13568 19499 13632
rect 19563 13568 19571 13632
rect 19251 12544 19571 13568
rect 19251 12480 19259 12544
rect 19323 12480 19339 12544
rect 19403 12480 19419 12544
rect 19483 12480 19499 12544
rect 19563 12480 19571 12544
rect 19251 11456 19571 12480
rect 19251 11392 19259 11456
rect 19323 11392 19339 11456
rect 19403 11392 19419 11456
rect 19483 11392 19499 11456
rect 19563 11392 19571 11456
rect 19251 10368 19571 11392
rect 19251 10304 19259 10368
rect 19323 10304 19339 10368
rect 19403 10304 19419 10368
rect 19483 10304 19499 10368
rect 19563 10304 19571 10368
rect 19251 9280 19571 10304
rect 19251 9216 19259 9280
rect 19323 9216 19339 9280
rect 19403 9216 19419 9280
rect 19483 9216 19499 9280
rect 19563 9216 19571 9280
rect 19251 8192 19571 9216
rect 19251 8128 19259 8192
rect 19323 8128 19339 8192
rect 19403 8128 19419 8192
rect 19483 8128 19499 8192
rect 19563 8128 19571 8192
rect 19251 7104 19571 8128
rect 19251 7040 19259 7104
rect 19323 7040 19339 7104
rect 19403 7040 19419 7104
rect 19483 7040 19499 7104
rect 19563 7040 19571 7104
rect 19251 6016 19571 7040
rect 19251 5952 19259 6016
rect 19323 5952 19339 6016
rect 19403 5952 19419 6016
rect 19483 5952 19499 6016
rect 19563 5952 19571 6016
rect 19251 4928 19571 5952
rect 19251 4864 19259 4928
rect 19323 4864 19339 4928
rect 19403 4864 19419 4928
rect 19483 4864 19499 4928
rect 19563 4864 19571 4928
rect 19251 3840 19571 4864
rect 19251 3776 19259 3840
rect 19323 3776 19339 3840
rect 19403 3776 19419 3840
rect 19483 3776 19499 3840
rect 19563 3776 19571 3840
rect 19251 2752 19571 3776
rect 19251 2688 19259 2752
rect 19323 2688 19339 2752
rect 19403 2688 19419 2752
rect 19483 2688 19499 2752
rect 19563 2688 19571 2752
rect 19251 1664 19571 2688
rect 19251 1600 19259 1664
rect 19323 1600 19339 1664
rect 19403 1600 19419 1664
rect 19483 1600 19499 1664
rect 19563 1600 19571 1664
rect 19251 576 19571 1600
rect 19251 512 19259 576
rect 19323 512 19339 576
rect 19403 512 19419 576
rect 19483 512 19499 576
rect 19563 512 19571 576
rect 19251 496 19571 512
use sky130_fd_sc_hd__inv_2  _03_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 17480 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _04_
timestamp 1693170804
transform 1 0 18124 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _05__10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 16560 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _05_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 16284 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_4  _06_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 18308 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 19136 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1693170804
transform -1 0 15456 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1693170804
transform 1 0 17296 0 -1 16864
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1693170804
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3220 0 1 544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_38
timestamp 1693170804
transform 1 0 4048 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_50
timestamp 1693170804
transform 1 0 5152 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 5796 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_61
timestamp 1693170804
transform 1 0 6164 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_65
timestamp 1693170804
transform 1 0 6532 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_77
timestamp 1693170804
transform 1 0 7636 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1693170804
transform 1 0 8188 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_85
timestamp 1693170804
transform 1 0 8372 0 1 544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_92
timestamp 1693170804
transform 1 0 9016 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_104 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 10120 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 10948 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_119
timestamp 1693170804
transform 1 0 11500 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_131
timestamp 1693170804
transform 1 0 12604 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1693170804
transform 1 0 13340 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_141 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 13524 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_146
timestamp 1693170804
transform 1 0 13984 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_158
timestamp 1693170804
transform 1 0 15088 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_166
timestamp 1693170804
transform 1 0 15824 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_169
timestamp 1693170804
transform 1 0 16100 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_173
timestamp 1693170804
transform 1 0 16468 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_185
timestamp 1693170804
transform 1 0 17572 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1693170804
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_200
timestamp 1693170804
transform 1 0 18952 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1693170804
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1693170804
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1693170804
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1693170804
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1693170804
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1693170804
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1693170804
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1693170804
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1693170804
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1693170804
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1693170804
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1693170804
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1693170804
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1693170804
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1693170804
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1693170804
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1693170804
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1693170804
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1693170804
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1693170804
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_193
timestamp 1693170804
transform 1 0 18308 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_201
timestamp 1693170804
transform 1 0 19044 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1693170804
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1693170804
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1693170804
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1693170804
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1693170804
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1693170804
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1693170804
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1693170804
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1693170804
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1693170804
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1693170804
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1693170804
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1693170804
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1693170804
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1693170804
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1693170804
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1693170804
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1693170804
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1693170804
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1693170804
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1693170804
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_197
timestamp 1693170804
transform 1 0 18676 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_201
timestamp 1693170804
transform 1 0 19044 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1693170804
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1693170804
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1693170804
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1693170804
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1693170804
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1693170804
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1693170804
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1693170804
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1693170804
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1693170804
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1693170804
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1693170804
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1693170804
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1693170804
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1693170804
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1693170804
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1693170804
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1693170804
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1693170804
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1693170804
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_193
timestamp 1693170804
transform 1 0 18308 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_201
timestamp 1693170804
transform 1 0 19044 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1693170804
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1693170804
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1693170804
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1693170804
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1693170804
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1693170804
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1693170804
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1693170804
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1693170804
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1693170804
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1693170804
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1693170804
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1693170804
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1693170804
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1693170804
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1693170804
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1693170804
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1693170804
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1693170804
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1693170804
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1693170804
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_197
timestamp 1693170804
transform 1 0 18676 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_201
timestamp 1693170804
transform 1 0 19044 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1693170804
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1693170804
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1693170804
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1693170804
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1693170804
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1693170804
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1693170804
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1693170804
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1693170804
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1693170804
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1693170804
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1693170804
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1693170804
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1693170804
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1693170804
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1693170804
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1693170804
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1693170804
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1693170804
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1693170804
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_193
timestamp 1693170804
transform 1 0 18308 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_201
timestamp 1693170804
transform 1 0 19044 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1693170804
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1693170804
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1693170804
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1693170804
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1693170804
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1693170804
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1693170804
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1693170804
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1693170804
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1693170804
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1693170804
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1693170804
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1693170804
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1693170804
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1693170804
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1693170804
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1693170804
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1693170804
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1693170804
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1693170804
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1693170804
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_197
timestamp 1693170804
transform 1 0 18676 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_201
timestamp 1693170804
transform 1 0 19044 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1693170804
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1693170804
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1693170804
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1693170804
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1693170804
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1693170804
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1693170804
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1693170804
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1693170804
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1693170804
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1693170804
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1693170804
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1693170804
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1693170804
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1693170804
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1693170804
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1693170804
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1693170804
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1693170804
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1693170804
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_193
timestamp 1693170804
transform 1 0 18308 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_201
timestamp 1693170804
transform 1 0 19044 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1693170804
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1693170804
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1693170804
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1693170804
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1693170804
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1693170804
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1693170804
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1693170804
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1693170804
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1693170804
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1693170804
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1693170804
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1693170804
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1693170804
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1693170804
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1693170804
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1693170804
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1693170804
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1693170804
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1693170804
transform 1 0 17940 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1693170804
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_197
timestamp 1693170804
transform 1 0 18676 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_201
timestamp 1693170804
transform 1 0 19044 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1693170804
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1693170804
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1693170804
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1693170804
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1693170804
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1693170804
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1693170804
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1693170804
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1693170804
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1693170804
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1693170804
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1693170804
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1693170804
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1693170804
transform 1 0 12052 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1693170804
transform 1 0 13156 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1693170804
transform 1 0 14260 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1693170804
transform 1 0 15364 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1693170804
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1693170804
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1693170804
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_193
timestamp 1693170804
transform 1 0 18308 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_201
timestamp 1693170804
transform 1 0 19044 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1693170804
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1693170804
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1693170804
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1693170804
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1693170804
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1693170804
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1693170804
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1693170804
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1693170804
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1693170804
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1693170804
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1693170804
transform 1 0 10580 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1693170804
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1693170804
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1693170804
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1693170804
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1693170804
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1693170804
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1693170804
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1693170804
transform 1 0 17940 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1693170804
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_197
timestamp 1693170804
transform 1 0 18676 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_201
timestamp 1693170804
transform 1 0 19044 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1693170804
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1693170804
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1693170804
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1693170804
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1693170804
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1693170804
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1693170804
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1693170804
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1693170804
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1693170804
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1693170804
transform 1 0 10212 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1693170804
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1693170804
transform 1 0 10948 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1693170804
transform 1 0 12052 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1693170804
transform 1 0 13156 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1693170804
transform 1 0 14260 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1693170804
transform 1 0 15364 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1693170804
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1693170804
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1693170804
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_193
timestamp 1693170804
transform 1 0 18308 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_201
timestamp 1693170804
transform 1 0 19044 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1693170804
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1693170804
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1693170804
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1693170804
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1693170804
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1693170804
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1693170804
transform 1 0 6532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1693170804
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1693170804
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1693170804
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1693170804
transform 1 0 9476 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1693170804
transform 1 0 10580 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1693170804
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1693170804
transform 1 0 12788 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1693170804
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1693170804
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1693170804
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1693170804
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1693170804
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1693170804
transform 1 0 17940 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1693170804
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_197
timestamp 1693170804
transform 1 0 18676 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_201
timestamp 1693170804
transform 1 0 19044 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1693170804
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1693170804
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1693170804
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1693170804
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1693170804
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1693170804
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1693170804
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1693170804
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1693170804
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1693170804
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1693170804
transform 1 0 10212 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1693170804
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1693170804
transform 1 0 10948 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1693170804
transform 1 0 12052 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1693170804
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1693170804
transform 1 0 14260 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1693170804
transform 1 0 15364 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1693170804
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1693170804
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1693170804
transform 1 0 17204 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_193
timestamp 1693170804
transform 1 0 18308 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_201
timestamp 1693170804
transform 1 0 19044 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1693170804
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1693170804
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1693170804
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1693170804
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1693170804
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1693170804
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1693170804
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1693170804
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1693170804
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1693170804
transform 1 0 8372 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1693170804
transform 1 0 9476 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1693170804
transform 1 0 10580 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1693170804
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1693170804
transform 1 0 12788 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1693170804
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1693170804
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1693170804
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1693170804
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1693170804
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1693170804
transform 1 0 17940 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1693170804
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_197
timestamp 1693170804
transform 1 0 18676 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_201
timestamp 1693170804
transform 1 0 19044 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1693170804
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1693170804
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1693170804
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1693170804
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1693170804
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1693170804
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1693170804
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1693170804
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1693170804
transform 1 0 8004 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1693170804
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1693170804
transform 1 0 10212 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1693170804
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1693170804
transform 1 0 10948 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1693170804
transform 1 0 12052 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1693170804
transform 1 0 13156 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1693170804
transform 1 0 14260 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1693170804
transform 1 0 15364 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1693170804
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1693170804
transform 1 0 16100 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1693170804
transform 1 0 17204 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_193
timestamp 1693170804
transform 1 0 18308 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_201
timestamp 1693170804
transform 1 0 19044 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1693170804
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1693170804
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1693170804
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1693170804
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1693170804
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1693170804
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1693170804
transform 1 0 6532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1693170804
transform 1 0 7636 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1693170804
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1693170804
transform 1 0 8372 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1693170804
transform 1 0 9476 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1693170804
transform 1 0 10580 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1693170804
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1693170804
transform 1 0 12788 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1693170804
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1693170804
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1693170804
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1693170804
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1693170804
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1693170804
transform 1 0 17940 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1693170804
transform 1 0 18492 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_197
timestamp 1693170804
transform 1 0 18676 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_201
timestamp 1693170804
transform 1 0 19044 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1693170804
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1693170804
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1693170804
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1693170804
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1693170804
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1693170804
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1693170804
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1693170804
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1693170804
transform 1 0 8004 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1693170804
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1693170804
transform 1 0 10212 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1693170804
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1693170804
transform 1 0 10948 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1693170804
transform 1 0 12052 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1693170804
transform 1 0 13156 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1693170804
transform 1 0 14260 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1693170804
transform 1 0 15364 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1693170804
transform 1 0 15916 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1693170804
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1693170804
transform 1 0 17204 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_193
timestamp 1693170804
transform 1 0 18308 0 -1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1693170804
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1693170804
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1693170804
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1693170804
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1693170804
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1693170804
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1693170804
transform 1 0 6532 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1693170804
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1693170804
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1693170804
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1693170804
transform 1 0 9476 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1693170804
transform 1 0 10580 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1693170804
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1693170804
transform 1 0 12788 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1693170804
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1693170804
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1693170804
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1693170804
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1693170804
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1693170804
transform 1 0 17940 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1693170804
transform 1 0 18492 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_197
timestamp 1693170804
transform 1 0 18676 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_201
timestamp 1693170804
transform 1 0 19044 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1693170804
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1693170804
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1693170804
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1693170804
transform 1 0 4140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1693170804
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1693170804
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1693170804
transform 1 0 5796 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1693170804
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1693170804
transform 1 0 8004 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1693170804
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1693170804
transform 1 0 10212 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1693170804
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1693170804
transform 1 0 10948 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1693170804
transform 1 0 12052 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1693170804
transform 1 0 13156 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1693170804
transform 1 0 14260 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1693170804
transform 1 0 15364 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1693170804
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1693170804
transform 1 0 16100 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1693170804
transform 1 0 17204 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_193
timestamp 1693170804
transform 1 0 18308 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_201
timestamp 1693170804
transform 1 0 19044 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1693170804
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1693170804
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1693170804
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1693170804
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1693170804
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1693170804
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1693170804
transform 1 0 6532 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1693170804
transform 1 0 7636 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1693170804
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1693170804
transform 1 0 8372 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1693170804
transform 1 0 9476 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1693170804
transform 1 0 10580 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1693170804
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1693170804
transform 1 0 12788 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1693170804
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1693170804
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1693170804
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1693170804
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1693170804
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1693170804
transform 1 0 17940 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1693170804
transform 1 0 18492 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_197
timestamp 1693170804
transform 1 0 18676 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_201
timestamp 1693170804
transform 1 0 19044 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1693170804
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1693170804
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1693170804
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1693170804
transform 1 0 4140 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1693170804
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1693170804
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1693170804
transform 1 0 5796 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1693170804
transform 1 0 6900 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1693170804
transform 1 0 8004 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1693170804
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1693170804
transform 1 0 10212 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1693170804
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1693170804
transform 1 0 10948 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1693170804
transform 1 0 12052 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1693170804
transform 1 0 13156 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1693170804
transform 1 0 14260 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1693170804
transform 1 0 15364 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1693170804
transform 1 0 15916 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1693170804
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1693170804
transform 1 0 17204 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_193
timestamp 1693170804
transform 1 0 18308 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_201
timestamp 1693170804
transform 1 0 19044 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1693170804
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1693170804
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1693170804
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1693170804
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1693170804
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1693170804
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1693170804
transform 1 0 6532 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1693170804
transform 1 0 7636 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1693170804
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1693170804
transform 1 0 8372 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1693170804
transform 1 0 9476 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1693170804
transform 1 0 10580 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1693170804
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1693170804
transform 1 0 12788 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1693170804
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1693170804
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1693170804
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1693170804
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1693170804
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1693170804
transform 1 0 17940 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1693170804
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_197
timestamp 1693170804
transform 1 0 18676 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_201
timestamp 1693170804
transform 1 0 19044 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1693170804
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1693170804
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1693170804
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1693170804
transform 1 0 4140 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1693170804
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1693170804
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1693170804
transform 1 0 5796 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1693170804
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1693170804
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1693170804
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1693170804
transform 1 0 10212 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1693170804
transform 1 0 10764 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1693170804
transform 1 0 10948 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1693170804
transform 1 0 12052 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1693170804
transform 1 0 13156 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1693170804
transform 1 0 14260 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1693170804
transform 1 0 15364 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1693170804
transform 1 0 15916 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1693170804
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1693170804
transform 1 0 17204 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_193
timestamp 1693170804
transform 1 0 18308 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_201
timestamp 1693170804
transform 1 0 19044 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1693170804
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1693170804
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1693170804
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1693170804
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1693170804
transform 1 0 4324 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1693170804
transform 1 0 5428 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1693170804
transform 1 0 6532 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1693170804
transform 1 0 7636 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1693170804
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1693170804
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1693170804
transform 1 0 9476 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1693170804
transform 1 0 10580 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1693170804
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1693170804
transform 1 0 12788 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1693170804
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1693170804
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1693170804
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1693170804
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1693170804
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1693170804
transform 1 0 17940 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1693170804
transform 1 0 18492 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_197
timestamp 1693170804
transform 1 0 18676 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_201
timestamp 1693170804
transform 1 0 19044 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1693170804
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1693170804
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1693170804
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1693170804
transform 1 0 4140 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1693170804
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1693170804
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1693170804
transform 1 0 5796 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1693170804
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1693170804
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1693170804
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1693170804
transform 1 0 10212 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1693170804
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1693170804
transform 1 0 10948 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1693170804
transform 1 0 12052 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1693170804
transform 1 0 13156 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1693170804
transform 1 0 14260 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1693170804
transform 1 0 15364 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1693170804
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1693170804
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1693170804
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_193
timestamp 1693170804
transform 1 0 18308 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_201
timestamp 1693170804
transform 1 0 19044 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1693170804
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1693170804
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1693170804
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1693170804
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1693170804
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1693170804
transform 1 0 5428 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1693170804
transform 1 0 6532 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1693170804
transform 1 0 7636 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1693170804
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1693170804
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1693170804
transform 1 0 9476 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1693170804
transform 1 0 10580 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1693170804
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1693170804
transform 1 0 12788 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1693170804
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1693170804
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1693170804
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1693170804
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1693170804
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1693170804
transform 1 0 17940 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1693170804
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_197
timestamp 1693170804
transform 1 0 18676 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_201
timestamp 1693170804
transform 1 0 19044 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1693170804
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1693170804
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1693170804
transform 1 0 3036 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1693170804
transform 1 0 4140 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1693170804
transform 1 0 5244 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1693170804
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1693170804
transform 1 0 5796 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1693170804
transform 1 0 6900 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1693170804
transform 1 0 8004 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1693170804
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1693170804
transform 1 0 10212 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1693170804
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1693170804
transform 1 0 10948 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1693170804
transform 1 0 12052 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1693170804
transform 1 0 13156 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1693170804
transform 1 0 14260 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1693170804
transform 1 0 15364 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1693170804
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1693170804
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1693170804
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_193
timestamp 1693170804
transform 1 0 18308 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_201
timestamp 1693170804
transform 1 0 19044 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1693170804
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1693170804
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1693170804
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1693170804
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1693170804
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1693170804
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1693170804
transform 1 0 6532 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1693170804
transform 1 0 7636 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1693170804
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1693170804
transform 1 0 8372 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1693170804
transform 1 0 9476 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1693170804
transform 1 0 10580 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1693170804
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1693170804
transform 1 0 12788 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1693170804
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1693170804
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1693170804
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1693170804
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1693170804
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1693170804
transform 1 0 17940 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1693170804
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_197
timestamp 1693170804
transform 1 0 18676 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_201
timestamp 1693170804
transform 1 0 19044 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1693170804
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1693170804
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1693170804
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1693170804
transform 1 0 4140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1693170804
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1693170804
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1693170804
transform 1 0 5796 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1693170804
transform 1 0 6900 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1693170804
transform 1 0 8004 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1693170804
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1693170804
transform 1 0 10212 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1693170804
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1693170804
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1693170804
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_137
timestamp 1693170804
transform 1 0 13156 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_141
timestamp 1693170804
transform 1 0 13524 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_162
timestamp 1693170804
transform 1 0 15456 0 -1 16864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1693170804
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_181
timestamp 1693170804
transform 1 0 17204 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1693170804
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1693170804
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1693170804
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1693170804
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1693170804
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1693170804
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1693170804
transform 1 0 6532 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1693170804
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1693170804
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1693170804
transform 1 0 8372 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1693170804
transform 1 0 9476 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1693170804
transform 1 0 10580 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1693170804
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1693170804
transform 1 0 12788 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1693170804
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1693170804
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1693170804
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_165
timestamp 1693170804
transform 1 0 15732 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_173
timestamp 1693170804
transform 1 0 16468 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_193
timestamp 1693170804
transform 1 0 18308 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_197
timestamp 1693170804
transform 1 0 18676 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_201
timestamp 1693170804
transform 1 0 19044 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1693170804
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1693170804
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1693170804
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1693170804
transform 1 0 4140 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1693170804
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1693170804
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1693170804
transform 1 0 5796 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1693170804
transform 1 0 6900 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1693170804
transform 1 0 8004 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1693170804
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1693170804
transform 1 0 10212 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1693170804
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1693170804
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1693170804
transform 1 0 12052 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1693170804
transform 1 0 13156 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1693170804
transform 1 0 14260 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1693170804
transform 1 0 15364 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1693170804
transform 1 0 15916 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1693170804
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_181
timestamp 1693170804
transform 1 0 17204 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1693170804
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1693170804
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1693170804
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1693170804
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1693170804
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1693170804
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1693170804
transform 1 0 6532 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1693170804
transform 1 0 7636 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1693170804
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1693170804
transform 1 0 8372 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1693170804
transform 1 0 9476 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1693170804
transform 1 0 10580 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1693170804
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1693170804
transform 1 0 12788 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1693170804
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1693170804
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1693170804
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_165
timestamp 1693170804
transform 1 0 15732 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_194
timestamp 1693170804
transform 1 0 18400 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_197
timestamp 1693170804
transform 1 0 18676 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_201
timestamp 1693170804
transform 1 0 19044 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1693170804
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1693170804
transform 1 0 1932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_27
timestamp 1693170804
transform 1 0 3036 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_29
timestamp 1693170804
transform 1 0 3220 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_41
timestamp 1693170804
transform 1 0 4324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1693170804
transform 1 0 5428 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1693170804
transform 1 0 5796 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1693170804
transform 1 0 6900 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_81
timestamp 1693170804
transform 1 0 8004 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_85
timestamp 1693170804
transform 1 0 8372 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_97
timestamp 1693170804
transform 1 0 9476 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1693170804
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1693170804
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1693170804
transform 1 0 12052 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_137
timestamp 1693170804
transform 1 0 13156 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_141
timestamp 1693170804
transform 1 0 13524 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_153
timestamp 1693170804
transform 1 0 14628 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1693170804
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_169
timestamp 1693170804
transform 1 0 16100 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_173
timestamp 1693170804
transform 1 0 16468 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_177
timestamp 1693170804
transform 1 0 16836 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_195
timestamp 1693170804
transform 1 0 18492 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_197
timestamp 1693170804
transform 1 0 18676 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_201
timestamp 1693170804
transform 1 0 19044 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 18492 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 17756 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp 1693170804
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1693170804
transform -1 0 19412 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp 1693170804
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1693170804
transform -1 0 19412 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp 1693170804
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1693170804
transform -1 0 19412 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp 1693170804
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1693170804
transform -1 0 19412 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp 1693170804
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1693170804
transform -1 0 19412 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp 1693170804
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1693170804
transform -1 0 19412 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp 1693170804
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1693170804
transform -1 0 19412 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp 1693170804
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1693170804
transform -1 0 19412 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp 1693170804
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1693170804
transform -1 0 19412 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp 1693170804
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1693170804
transform -1 0 19412 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp 1693170804
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1693170804
transform -1 0 19412 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp 1693170804
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1693170804
transform -1 0 19412 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp 1693170804
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1693170804
transform -1 0 19412 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp 1693170804
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1693170804
transform -1 0 19412 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp 1693170804
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1693170804
transform -1 0 19412 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp 1693170804
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1693170804
transform -1 0 19412 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp 1693170804
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1693170804
transform -1 0 19412 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp 1693170804
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1693170804
transform -1 0 19412 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp 1693170804
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1693170804
transform -1 0 19412 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp 1693170804
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1693170804
transform -1 0 19412 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp 1693170804
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1693170804
transform -1 0 19412 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp 1693170804
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1693170804
transform -1 0 19412 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp 1693170804
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1693170804
transform -1 0 19412 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp 1693170804
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1693170804
transform -1 0 19412 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp 1693170804
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1693170804
transform -1 0 19412 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp 1693170804
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1693170804
transform -1 0 19412 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp 1693170804
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1693170804
transform -1 0 19412 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp 1693170804
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1693170804
transform -1 0 19412 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp 1693170804
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1693170804
transform -1 0 19412 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp 1693170804
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1693170804
transform -1 0 19412 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp 1693170804
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1693170804
transform -1 0 19412 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp 1693170804
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1693170804
transform -1 0 19412 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp 1693170804
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1693170804
transform -1 0 19412 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp 1693170804
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1693170804
transform -1 0 19412 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  r2r_dac_control_2
timestamp 1693170804
transform 1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  r2r_dac_control_3
timestamp 1693170804
transform -1 0 4048 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  r2r_dac_control_4
timestamp 1693170804
transform -1 0 6532 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  r2r_dac_control_5
timestamp 1693170804
transform -1 0 9016 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  r2r_dac_control_6
timestamp 1693170804
transform -1 0 11500 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  r2r_dac_control_7
timestamp 1693170804
transform -1 0 13984 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  r2r_dac_control_8
timestamp 1693170804
transform -1 0 16468 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  r2r_dac_control_9
timestamp 1693170804
transform -1 0 18952 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 1693170804
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 1693170804
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1693170804
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1693170804
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1693170804
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1693170804
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_75
timestamp 1693170804
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_76
timestamp 1693170804
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_77
timestamp 1693170804
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_78
timestamp 1693170804
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_79
timestamp 1693170804
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_80
timestamp 1693170804
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_81
timestamp 1693170804
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_82
timestamp 1693170804
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_83
timestamp 1693170804
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_84
timestamp 1693170804
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_85
timestamp 1693170804
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_86
timestamp 1693170804
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_87
timestamp 1693170804
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_88
timestamp 1693170804
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_89
timestamp 1693170804
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_90
timestamp 1693170804
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_91
timestamp 1693170804
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_92
timestamp 1693170804
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_93
timestamp 1693170804
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_94
timestamp 1693170804
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_95
timestamp 1693170804
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_96
timestamp 1693170804
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_97
timestamp 1693170804
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_98
timestamp 1693170804
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_99
timestamp 1693170804
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_100
timestamp 1693170804
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_101
timestamp 1693170804
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_102
timestamp 1693170804
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_103
timestamp 1693170804
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_104
timestamp 1693170804
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_105
timestamp 1693170804
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp 1693170804
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp 1693170804
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_108
timestamp 1693170804
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_109
timestamp 1693170804
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp 1693170804
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp 1693170804
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp 1693170804
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_113
timestamp 1693170804
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_114
timestamp 1693170804
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_115
timestamp 1693170804
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_116
timestamp 1693170804
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_117
timestamp 1693170804
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_118
timestamp 1693170804
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_119
timestamp 1693170804
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_120
timestamp 1693170804
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_121
timestamp 1693170804
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_122
timestamp 1693170804
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_123
timestamp 1693170804
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_124
timestamp 1693170804
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_125
timestamp 1693170804
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_126
timestamp 1693170804
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_127
timestamp 1693170804
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_128
timestamp 1693170804
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_129
timestamp 1693170804
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_130
timestamp 1693170804
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_131
timestamp 1693170804
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_132
timestamp 1693170804
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_133
timestamp 1693170804
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_134
timestamp 1693170804
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_135
timestamp 1693170804
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_136
timestamp 1693170804
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_137
timestamp 1693170804
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_138
timestamp 1693170804
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_139
timestamp 1693170804
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_140
timestamp 1693170804
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_141
timestamp 1693170804
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_142
timestamp 1693170804
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_143
timestamp 1693170804
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_144
timestamp 1693170804
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_145
timestamp 1693170804
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_146
timestamp 1693170804
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_147
timestamp 1693170804
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_148
timestamp 1693170804
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_149
timestamp 1693170804
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_150
timestamp 1693170804
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_151
timestamp 1693170804
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_152
timestamp 1693170804
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_153
timestamp 1693170804
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_154
timestamp 1693170804
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_155
timestamp 1693170804
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_156
timestamp 1693170804
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_157
timestamp 1693170804
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_158
timestamp 1693170804
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_159
timestamp 1693170804
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_160
timestamp 1693170804
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_161
timestamp 1693170804
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_162
timestamp 1693170804
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_163
timestamp 1693170804
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_164
timestamp 1693170804
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_165
timestamp 1693170804
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_166
timestamp 1693170804
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_167
timestamp 1693170804
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_168
timestamp 1693170804
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_169
timestamp 1693170804
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_170
timestamp 1693170804
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_171
timestamp 1693170804
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_172
timestamp 1693170804
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_173
timestamp 1693170804
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_174
timestamp 1693170804
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_175
timestamp 1693170804
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_176
timestamp 1693170804
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_177
timestamp 1693170804
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_178
timestamp 1693170804
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_179
timestamp 1693170804
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_180
timestamp 1693170804
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_181
timestamp 1693170804
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_182
timestamp 1693170804
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_183
timestamp 1693170804
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_184
timestamp 1693170804
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_185
timestamp 1693170804
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_186
timestamp 1693170804
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_187
timestamp 1693170804
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_188
timestamp 1693170804
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_189
timestamp 1693170804
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_190
timestamp 1693170804
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_191
timestamp 1693170804
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_192
timestamp 1693170804
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_193
timestamp 1693170804
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
<< labels >>
flabel metal4 s 5106 496 5426 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 9821 496 10141 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 14536 496 14856 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 19251 496 19571 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2749 496 3069 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7464 496 7784 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12179 496 12499 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 16894 496 17214 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 19062 19600 19118 20000 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal3 s 19600 9800 20000 9920 0 FreeSans 480 0 0 0 cnt_zero
port 3 nsew signal tristate
flabel metal2 s 15750 19600 15806 20000 0 FreeSans 224 90 0 0 data[0]
port 4 nsew signal input
flabel metal2 s 14094 19600 14150 20000 0 FreeSans 224 90 0 0 data[1]
port 5 nsew signal input
flabel metal2 s 12438 19600 12494 20000 0 FreeSans 224 90 0 0 data[2]
port 6 nsew signal input
flabel metal2 s 10782 19600 10838 20000 0 FreeSans 224 90 0 0 data[3]
port 7 nsew signal input
flabel metal2 s 9126 19600 9182 20000 0 FreeSans 224 90 0 0 data[4]
port 8 nsew signal input
flabel metal2 s 7470 19600 7526 20000 0 FreeSans 224 90 0 0 data[5]
port 9 nsew signal input
flabel metal2 s 5814 19600 5870 20000 0 FreeSans 224 90 0 0 data[6]
port 10 nsew signal input
flabel metal2 s 4158 19600 4214 20000 0 FreeSans 224 90 0 0 data[7]
port 11 nsew signal input
flabel metal2 s 2502 19600 2558 20000 0 FreeSans 224 90 0 0 ext_data
port 12 nsew signal input
flabel metal2 s 846 19600 902 20000 0 FreeSans 224 90 0 0 load_divider
port 13 nsew signal input
flabel metal2 s 17406 19600 17462 20000 0 FreeSans 224 90 0 0 n_rst
port 14 nsew signal input
flabel metal2 s 1214 0 1270 400 0 FreeSans 224 90 0 0 r2r_out[0]
port 15 nsew signal tristate
flabel metal2 s 3698 0 3754 400 0 FreeSans 224 90 0 0 r2r_out[1]
port 16 nsew signal tristate
flabel metal2 s 6182 0 6238 400 0 FreeSans 224 90 0 0 r2r_out[2]
port 17 nsew signal tristate
flabel metal2 s 8666 0 8722 400 0 FreeSans 224 90 0 0 r2r_out[3]
port 18 nsew signal tristate
flabel metal2 s 11150 0 11206 400 0 FreeSans 224 90 0 0 r2r_out[4]
port 19 nsew signal tristate
flabel metal2 s 13634 0 13690 400 0 FreeSans 224 90 0 0 r2r_out[5]
port 20 nsew signal tristate
flabel metal2 s 16118 0 16174 400 0 FreeSans 224 90 0 0 r2r_out[6]
port 21 nsew signal tristate
flabel metal2 s 18602 0 18658 400 0 FreeSans 224 90 0 0 r2r_out[7]
port 22 nsew signal tristate
rlabel via1 10061 19040 10061 19040 0 VGND
rlabel metal1 9982 18496 9982 18496 0 VPWR
rlabel metal1 17664 17170 17664 17170 0 _00_
rlabel metal1 18039 18122 18039 18122 0 _01_
rlabel metal2 19090 18710 19090 18710 0 clk
rlabel metal1 17480 16694 17480 16694 0 clknet_0_clk
rlabel metal1 15226 18190 15226 18190 0 clknet_1_0__leaf_clk
rlabel metal1 18446 17102 18446 17102 0 clknet_1_1__leaf_clk
rlabel metal1 17526 18836 17526 18836 0 n_rst
rlabel metal1 18170 18224 18170 18224 0 net1
rlabel metal2 16606 18496 16606 18496 0 net10
rlabel metal1 17434 18768 17434 18768 0 net11
rlabel metal3 19420 9860 19420 9860 0 net2
rlabel metal2 3726 415 3726 415 0 net3
rlabel metal2 6210 415 6210 415 0 net4
rlabel metal2 8694 415 8694 415 0 net5
rlabel metal2 11178 415 11178 415 0 net6
rlabel metal2 13662 415 13662 415 0 net7
rlabel metal2 16146 415 16146 415 0 net8
rlabel metal2 18630 415 18630 415 0 net9
rlabel metal2 1242 8796 1242 8796 0 r2r_out[0]
rlabel metal1 18216 18394 18216 18394 0 rst
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
