magic
tech sky130A
magscale 1 2
timestamp 1720441783
<< error_p >>
rect -29 117 29 123
rect -29 83 -17 117
rect -29 77 29 83
rect -29 -83 29 -77
rect -29 -117 -17 -83
rect -29 -123 29 -117
<< nmos >>
rect -30 -45 30 45
<< ndiff >>
rect -88 33 -30 45
rect -88 -33 -76 33
rect -42 -33 -30 33
rect -88 -45 -30 -33
rect 30 33 88 45
rect 30 -33 42 33
rect 76 -33 88 33
rect 30 -45 88 -33
<< ndiffc >>
rect -76 -33 -42 33
rect 42 -33 76 33
<< poly >>
rect -33 117 33 133
rect -33 83 -17 117
rect 17 83 33 117
rect -33 67 33 83
rect -30 45 30 67
rect -30 -67 30 -45
rect -33 -83 33 -67
rect -33 -117 -17 -83
rect 17 -117 33 -83
rect -33 -133 33 -117
<< polycont >>
rect -17 83 17 117
rect -17 -117 17 -83
<< locali >>
rect -33 83 -17 117
rect 17 83 33 117
rect -76 33 -42 49
rect -76 -49 -42 -33
rect 42 33 76 49
rect 42 -49 76 -33
rect -33 -117 -17 -83
rect 17 -117 33 -83
<< viali >>
rect -17 83 17 117
rect -76 -33 -42 33
rect 42 -33 76 33
rect -17 -117 17 -83
<< metal1 >>
rect -29 117 29 123
rect -29 83 -17 117
rect 17 83 29 117
rect -29 77 29 83
rect -82 33 -36 45
rect -82 -33 -76 33
rect -42 -33 -36 33
rect -82 -45 -36 -33
rect 36 33 82 45
rect 36 -33 42 33
rect 76 -33 82 33
rect 36 -45 82 -33
rect -29 -83 29 -77
rect -29 -117 -17 -83
rect 17 -117 29 -83
rect -29 -123 29 -117
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.450 l 0.300 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
