magic
tech sky130A
timestamp 1725627062
<< pwell >>
rect -139 -529 139 529
<< mvnmos >>
rect -25 -400 25 400
<< mvndiff >>
rect -54 394 -25 400
rect -54 -394 -48 394
rect -31 -394 -25 394
rect -54 -400 -25 -394
rect 25 394 54 400
rect 25 -394 31 394
rect 48 -394 54 394
rect 25 -400 54 -394
<< mvndiffc >>
rect -48 -394 -31 394
rect 31 -394 48 394
<< mvpsubdiff >>
rect -121 505 121 511
rect -121 488 -67 505
rect 67 488 121 505
rect -121 482 121 488
rect -121 457 -92 482
rect -121 -457 -115 457
rect -98 -457 -92 457
rect 92 457 121 482
rect -121 -482 -92 -457
rect 92 -457 98 457
rect 115 -457 121 457
rect 92 -482 121 -457
rect -121 -488 121 -482
rect -121 -505 -67 -488
rect 67 -505 121 -488
rect -121 -511 121 -505
<< mvpsubdiffcont >>
rect -67 488 67 505
rect -115 -457 -98 457
rect 98 -457 115 457
rect -67 -505 67 -488
<< poly >>
rect -25 436 25 444
rect -25 419 -17 436
rect 17 419 25 436
rect -25 400 25 419
rect -25 -419 25 -400
rect -25 -436 -17 -419
rect 17 -436 25 -419
rect -25 -444 25 -436
<< polycont >>
rect -17 419 17 436
rect -17 -436 17 -419
<< locali >>
rect -115 488 -67 505
rect 67 488 115 505
rect -115 457 -98 488
rect 98 457 115 488
rect -25 419 -17 436
rect 17 419 25 436
rect -48 394 -31 402
rect -48 -402 -31 -394
rect 31 394 48 402
rect 31 -402 48 -394
rect -25 -436 -17 -419
rect 17 -436 25 -419
rect -115 -488 -98 -457
rect 98 -488 115 -457
rect -115 -505 -67 -488
rect 67 -505 115 -488
<< viali >>
rect -17 419 17 436
rect -48 -394 -31 394
rect 31 -394 48 394
rect -17 -436 17 -419
<< metal1 >>
rect -23 436 23 439
rect -23 419 -17 436
rect 17 419 23 436
rect -23 416 23 419
rect -51 394 -28 400
rect -51 -394 -48 394
rect -31 -394 -28 394
rect -51 -400 -28 -394
rect 28 394 51 400
rect 28 -394 31 394
rect 48 -394 51 394
rect 28 -400 51 -394
rect -23 -419 23 -416
rect -23 -436 -17 -419
rect 17 -436 23 -419
rect -23 -439 23 -436
<< properties >>
string FIXED_BBOX -106 -496 106 496
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 8 l 0.50 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__nfet_g5v0d10v5_F263WR gencell
<< end >>
