magic
tech sky130A
magscale 1 2
timestamp 1725626266
<< metal3 >>
rect -8298 5172 -2926 5200
rect -8298 148 -3010 5172
rect -2946 148 -2926 5172
rect -8298 120 -2926 148
rect -2686 5172 2686 5200
rect -2686 148 2602 5172
rect 2666 148 2686 5172
rect -2686 120 2686 148
rect 2926 5172 8298 5200
rect 2926 148 8214 5172
rect 8278 148 8298 5172
rect 2926 120 8298 148
rect -8298 -148 -2926 -120
rect -8298 -5172 -3010 -148
rect -2946 -5172 -2926 -148
rect -8298 -5200 -2926 -5172
rect -2686 -148 2686 -120
rect -2686 -5172 2602 -148
rect 2666 -5172 2686 -148
rect -2686 -5200 2686 -5172
rect 2926 -148 8298 -120
rect 2926 -5172 8214 -148
rect 8278 -5172 8298 -148
rect 2926 -5200 8298 -5172
<< via3 >>
rect -3010 148 -2946 5172
rect 2602 148 2666 5172
rect 8214 148 8278 5172
rect -3010 -5172 -2946 -148
rect 2602 -5172 2666 -148
rect 8214 -5172 8278 -148
<< mimcap >>
rect -8258 5120 -3258 5160
rect -8258 200 -8218 5120
rect -3298 200 -3258 5120
rect -8258 160 -3258 200
rect -2646 5120 2354 5160
rect -2646 200 -2606 5120
rect 2314 200 2354 5120
rect -2646 160 2354 200
rect 2966 5120 7966 5160
rect 2966 200 3006 5120
rect 7926 200 7966 5120
rect 2966 160 7966 200
rect -8258 -200 -3258 -160
rect -8258 -5120 -8218 -200
rect -3298 -5120 -3258 -200
rect -8258 -5160 -3258 -5120
rect -2646 -200 2354 -160
rect -2646 -5120 -2606 -200
rect 2314 -5120 2354 -200
rect -2646 -5160 2354 -5120
rect 2966 -200 7966 -160
rect 2966 -5120 3006 -200
rect 7926 -5120 7966 -200
rect 2966 -5160 7966 -5120
<< mimcapcontact >>
rect -8218 200 -3298 5120
rect -2606 200 2314 5120
rect 3006 200 7926 5120
rect -8218 -5120 -3298 -200
rect -2606 -5120 2314 -200
rect 3006 -5120 7926 -200
<< metal4 >>
rect -5810 5121 -5706 5320
rect -3030 5172 -2926 5320
rect -8219 5120 -3297 5121
rect -8219 200 -8218 5120
rect -3298 200 -3297 5120
rect -8219 199 -3297 200
rect -5810 -199 -5706 199
rect -3030 148 -3010 5172
rect -2946 148 -2926 5172
rect -198 5121 -94 5320
rect 2582 5172 2686 5320
rect -2607 5120 2315 5121
rect -2607 200 -2606 5120
rect 2314 200 2315 5120
rect -2607 199 2315 200
rect -3030 -148 -2926 148
rect -8219 -200 -3297 -199
rect -8219 -5120 -8218 -200
rect -3298 -5120 -3297 -200
rect -8219 -5121 -3297 -5120
rect -5810 -5320 -5706 -5121
rect -3030 -5172 -3010 -148
rect -2946 -5172 -2926 -148
rect -198 -199 -94 199
rect 2582 148 2602 5172
rect 2666 148 2686 5172
rect 5414 5121 5518 5320
rect 8194 5172 8298 5320
rect 3005 5120 7927 5121
rect 3005 200 3006 5120
rect 7926 200 7927 5120
rect 3005 199 7927 200
rect 2582 -148 2686 148
rect -2607 -200 2315 -199
rect -2607 -5120 -2606 -200
rect 2314 -5120 2315 -200
rect -2607 -5121 2315 -5120
rect -3030 -5320 -2926 -5172
rect -198 -5320 -94 -5121
rect 2582 -5172 2602 -148
rect 2666 -5172 2686 -148
rect 5414 -199 5518 199
rect 8194 148 8214 5172
rect 8278 148 8298 5172
rect 8194 -148 8298 148
rect 3005 -200 7927 -199
rect 3005 -5120 3006 -200
rect 7926 -5120 7927 -200
rect 3005 -5121 7927 -5120
rect 2582 -5320 2686 -5172
rect 5414 -5320 5518 -5121
rect 8194 -5172 8214 -148
rect 8278 -5172 8298 -148
rect 8194 -5320 8298 -5172
<< properties >>
string FIXED_BBOX 2926 120 8006 5200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25.00 l 25 val 1.269k carea 2.00 cperi 0.19 nx 3 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string sky130_fd_pr__cap_mim_m3_1_WFMHFS parameters
<< end >>
