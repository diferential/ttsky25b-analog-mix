magic
tech sky130A
magscale 1 2
timestamp 1762739948
<< metal3 >>
rect -386 212 386 240
rect -386 -212 302 212
rect 366 -212 386 212
rect -386 -240 386 -212
<< via3 >>
rect 302 -212 366 212
<< mimcap >>
rect -346 160 54 200
rect -346 -160 -306 160
rect 14 -160 54 160
rect -346 -200 54 -160
<< mimcapcontact >>
rect -306 -160 14 160
<< metal4 >>
rect 286 212 382 228
rect -307 160 15 161
rect -307 -160 -306 160
rect 14 -160 15 160
rect -307 -161 15 -160
rect 286 -212 302 212
rect 366 -212 382 212
rect 286 -228 382 -212
<< properties >>
string FIXED_BBOX -386 -240 94 240
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string sky130_fd_pr__cap_mim_m3_1_FJFAMD parameters
<< end >>
