magic
tech sky130A
magscale 1 2
timestamp 1720618976
<< nwell >>
rect -193 -112 193 112
<< pmoslvt >>
rect -99 -50 -29 50
rect 29 -50 99 50
<< pdiff >>
rect -157 38 -99 50
rect -157 -38 -145 38
rect -111 -38 -99 38
rect -157 -50 -99 -38
rect -29 38 29 50
rect -29 -38 -17 38
rect 17 -38 29 38
rect -29 -50 29 -38
rect 99 38 157 50
rect 99 -38 111 38
rect 145 -38 157 38
rect 99 -50 157 -38
<< pdiffc >>
rect -145 -38 -111 38
rect -17 -38 17 38
rect 111 -38 145 38
<< poly >>
rect -99 50 -29 76
rect 29 50 99 76
rect -99 -76 -29 -50
rect 29 -76 99 -50
<< locali >>
rect -145 38 -111 54
rect -145 -54 -111 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 111 38 145 54
rect 111 -54 145 -38
<< viali >>
rect -145 -38 -111 38
rect -17 -38 17 38
rect 111 -38 145 38
<< metal1 >>
rect -151 38 -105 50
rect -151 -38 -145 38
rect -111 -38 -105 38
rect -151 -50 -105 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 105 38 151 50
rect 105 -38 111 38
rect 145 -38 151 38
rect 105 -50 151 -38
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 0.5 l 0.35 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
