magic
tech sky130A
magscale 1 2
timestamp 1718373125
<< pwell >>
rect -647 -403 647 403
<< nmos >>
rect -447 109 -417 193
rect -351 109 -321 193
rect -255 109 -225 193
rect -159 109 -129 193
rect -63 109 -33 193
rect 33 109 63 193
rect 129 109 159 193
rect 225 109 255 193
rect 321 109 351 193
rect 417 109 447 193
rect -447 -193 -417 -109
rect -351 -193 -321 -109
rect -255 -193 -225 -109
rect -159 -193 -129 -109
rect -63 -193 -33 -109
rect 33 -193 63 -109
rect 129 -193 159 -109
rect 225 -193 255 -109
rect 321 -193 351 -109
rect 417 -193 447 -109
<< ndiff >>
rect -509 181 -447 193
rect -509 121 -497 181
rect -463 121 -447 181
rect -509 109 -447 121
rect -417 181 -351 193
rect -417 121 -401 181
rect -367 121 -351 181
rect -417 109 -351 121
rect -321 181 -255 193
rect -321 121 -305 181
rect -271 121 -255 181
rect -321 109 -255 121
rect -225 181 -159 193
rect -225 121 -209 181
rect -175 121 -159 181
rect -225 109 -159 121
rect -129 181 -63 193
rect -129 121 -113 181
rect -79 121 -63 181
rect -129 109 -63 121
rect -33 181 33 193
rect -33 121 -17 181
rect 17 121 33 181
rect -33 109 33 121
rect 63 181 129 193
rect 63 121 79 181
rect 113 121 129 181
rect 63 109 129 121
rect 159 181 225 193
rect 159 121 175 181
rect 209 121 225 181
rect 159 109 225 121
rect 255 181 321 193
rect 255 121 271 181
rect 305 121 321 181
rect 255 109 321 121
rect 351 181 417 193
rect 351 121 367 181
rect 401 121 417 181
rect 351 109 417 121
rect 447 181 509 193
rect 447 121 463 181
rect 497 121 509 181
rect 447 109 509 121
rect -509 -121 -447 -109
rect -509 -181 -497 -121
rect -463 -181 -447 -121
rect -509 -193 -447 -181
rect -417 -121 -351 -109
rect -417 -181 -401 -121
rect -367 -181 -351 -121
rect -417 -193 -351 -181
rect -321 -121 -255 -109
rect -321 -181 -305 -121
rect -271 -181 -255 -121
rect -321 -193 -255 -181
rect -225 -121 -159 -109
rect -225 -181 -209 -121
rect -175 -181 -159 -121
rect -225 -193 -159 -181
rect -129 -121 -63 -109
rect -129 -181 -113 -121
rect -79 -181 -63 -121
rect -129 -193 -63 -181
rect -33 -121 33 -109
rect -33 -181 -17 -121
rect 17 -181 33 -121
rect -33 -193 33 -181
rect 63 -121 129 -109
rect 63 -181 79 -121
rect 113 -181 129 -121
rect 63 -193 129 -181
rect 159 -121 225 -109
rect 159 -181 175 -121
rect 209 -181 225 -121
rect 159 -193 225 -181
rect 255 -121 321 -109
rect 255 -181 271 -121
rect 305 -181 321 -121
rect 255 -193 321 -181
rect 351 -121 417 -109
rect 351 -181 367 -121
rect 401 -181 417 -121
rect 351 -193 417 -181
rect 447 -121 509 -109
rect 447 -181 463 -121
rect 497 -181 509 -121
rect 447 -193 509 -181
<< ndiffc >>
rect -497 121 -463 181
rect -401 121 -367 181
rect -305 121 -271 181
rect -209 121 -175 181
rect -113 121 -79 181
rect -17 121 17 181
rect 79 121 113 181
rect 175 121 209 181
rect 271 121 305 181
rect 367 121 401 181
rect 463 121 497 181
rect -497 -181 -463 -121
rect -401 -181 -367 -121
rect -305 -181 -271 -121
rect -209 -181 -175 -121
rect -113 -181 -79 -121
rect -17 -181 17 -121
rect 79 -181 113 -121
rect 175 -181 209 -121
rect 271 -181 305 -121
rect 367 -181 401 -121
rect 463 -181 497 -121
<< psubdiff >>
rect -611 333 -515 367
rect 515 333 611 367
rect -611 271 -577 333
rect 577 271 611 333
rect -611 -333 -577 -271
rect 577 -333 611 -271
rect -611 -367 -515 -333
rect 515 -367 611 -333
<< psubdiffcont >>
rect -515 333 515 367
rect -611 -271 -577 271
rect 577 -271 611 271
rect -515 -367 515 -333
<< poly >>
rect -465 265 -399 281
rect -465 231 -449 265
rect -415 231 -399 265
rect -465 215 -399 231
rect -273 265 -207 281
rect -273 231 -257 265
rect -223 231 -207 265
rect -447 193 -417 215
rect -351 193 -321 219
rect -273 215 -207 231
rect -81 265 -15 281
rect -81 231 -65 265
rect -31 231 -15 265
rect -255 193 -225 215
rect -159 193 -129 219
rect -81 215 -15 231
rect 111 265 177 281
rect 111 231 127 265
rect 161 231 177 265
rect -63 193 -33 215
rect 33 193 63 219
rect 111 215 177 231
rect 303 265 369 281
rect 303 231 319 265
rect 353 231 369 265
rect 129 193 159 215
rect 225 193 255 219
rect 303 215 369 231
rect 321 193 351 215
rect 417 193 447 219
rect -447 83 -417 109
rect -351 87 -321 109
rect -369 71 -303 87
rect -255 83 -225 109
rect -159 87 -129 109
rect -369 37 -353 71
rect -319 37 -303 71
rect -369 21 -303 37
rect -177 71 -111 87
rect -63 83 -33 109
rect 33 87 63 109
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 129 83 159 109
rect 225 87 255 109
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 207 71 273 87
rect 321 83 351 109
rect 417 87 447 109
rect 207 37 223 71
rect 257 37 273 71
rect 207 21 273 37
rect 399 71 465 87
rect 399 37 415 71
rect 449 37 465 71
rect 399 21 465 37
rect -369 -37 -303 -21
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -447 -109 -417 -83
rect -369 -87 -303 -71
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -351 -109 -321 -87
rect -255 -109 -225 -83
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -159 -109 -129 -87
rect -63 -109 -33 -83
rect 15 -87 81 -71
rect 207 -37 273 -21
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 33 -109 63 -87
rect 129 -109 159 -83
rect 207 -87 273 -71
rect 399 -37 465 -21
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 225 -109 255 -87
rect 321 -109 351 -83
rect 399 -87 465 -71
rect 417 -109 447 -87
rect -447 -215 -417 -193
rect -465 -231 -399 -215
rect -351 -219 -321 -193
rect -255 -215 -225 -193
rect -465 -265 -449 -231
rect -415 -265 -399 -231
rect -465 -281 -399 -265
rect -273 -231 -207 -215
rect -159 -219 -129 -193
rect -63 -215 -33 -193
rect -273 -265 -257 -231
rect -223 -265 -207 -231
rect -273 -281 -207 -265
rect -81 -231 -15 -215
rect 33 -219 63 -193
rect 129 -215 159 -193
rect -81 -265 -65 -231
rect -31 -265 -15 -231
rect -81 -281 -15 -265
rect 111 -231 177 -215
rect 225 -219 255 -193
rect 321 -215 351 -193
rect 111 -265 127 -231
rect 161 -265 177 -231
rect 111 -281 177 -265
rect 303 -231 369 -215
rect 417 -219 447 -193
rect 303 -265 319 -231
rect 353 -265 369 -231
rect 303 -281 369 -265
<< polycont >>
rect -449 231 -415 265
rect -257 231 -223 265
rect -65 231 -31 265
rect 127 231 161 265
rect 319 231 353 265
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect -449 -265 -415 -231
rect -257 -265 -223 -231
rect -65 -265 -31 -231
rect 127 -265 161 -231
rect 319 -265 353 -231
<< locali >>
rect -611 333 -515 367
rect 515 333 611 367
rect -611 271 -577 333
rect 577 271 611 333
rect -465 231 -449 265
rect -415 231 -399 265
rect -273 231 -257 265
rect -223 231 -207 265
rect -81 231 -65 265
rect -31 231 -15 265
rect 111 231 127 265
rect 161 231 177 265
rect 303 231 319 265
rect 353 231 369 265
rect -497 181 -463 197
rect -497 105 -463 121
rect -401 181 -367 197
rect -401 105 -367 121
rect -305 181 -271 197
rect -305 105 -271 121
rect -209 181 -175 197
rect -209 105 -175 121
rect -113 181 -79 197
rect -113 105 -79 121
rect -17 181 17 197
rect -17 105 17 121
rect 79 181 113 197
rect 79 105 113 121
rect 175 181 209 197
rect 175 105 209 121
rect 271 181 305 197
rect 271 105 305 121
rect 367 181 401 197
rect 367 105 401 121
rect 463 181 497 197
rect 463 105 497 121
rect -369 37 -353 71
rect -319 37 -303 71
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect 207 37 223 71
rect 257 37 273 71
rect 399 37 415 71
rect 449 37 465 71
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 399 -71 415 -37
rect 449 -71 465 -37
rect -497 -121 -463 -105
rect -497 -197 -463 -181
rect -401 -121 -367 -105
rect -401 -197 -367 -181
rect -305 -121 -271 -105
rect -305 -197 -271 -181
rect -209 -121 -175 -105
rect -209 -197 -175 -181
rect -113 -121 -79 -105
rect -113 -197 -79 -181
rect -17 -121 17 -105
rect -17 -197 17 -181
rect 79 -121 113 -105
rect 79 -197 113 -181
rect 175 -121 209 -105
rect 175 -197 209 -181
rect 271 -121 305 -105
rect 271 -197 305 -181
rect 367 -121 401 -105
rect 367 -197 401 -181
rect 463 -121 497 -105
rect 463 -197 497 -181
rect -465 -265 -449 -231
rect -415 -265 -399 -231
rect -273 -265 -257 -231
rect -223 -265 -207 -231
rect -81 -265 -65 -231
rect -31 -265 -15 -231
rect 111 -265 127 -231
rect 161 -265 177 -231
rect 303 -265 319 -231
rect 353 -265 369 -231
rect -611 -333 -577 -271
rect 577 -333 611 -271
rect -611 -367 -515 -333
rect 515 -367 611 -333
<< properties >>
string FIXED_BBOX -594 -350 594 350
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.150 m 2 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
