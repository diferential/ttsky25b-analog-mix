magic
tech sky130A
magscale 1 2
timestamp 1762739948
<< pwell >>
rect -515 -327 515 327
<< mvnmos >>
rect -287 -131 -187 69
rect -129 -131 -29 69
rect 29 -131 129 69
rect 187 -131 287 69
<< mvndiff >>
rect -345 57 -287 69
rect -345 -119 -333 57
rect -299 -119 -287 57
rect -345 -131 -287 -119
rect -187 57 -129 69
rect -187 -119 -175 57
rect -141 -119 -129 57
rect -187 -131 -129 -119
rect -29 57 29 69
rect -29 -119 -17 57
rect 17 -119 29 57
rect -29 -131 29 -119
rect 129 57 187 69
rect 129 -119 141 57
rect 175 -119 187 57
rect 129 -131 187 -119
rect 287 57 345 69
rect 287 -119 299 57
rect 333 -119 345 57
rect 287 -131 345 -119
<< mvndiffc >>
rect -333 -119 -299 57
rect -175 -119 -141 57
rect -17 -119 17 57
rect 141 -119 175 57
rect 299 -119 333 57
<< mvpsubdiff >>
rect -479 279 479 291
rect -479 245 -371 279
rect 371 245 479 279
rect -479 233 479 245
rect -479 183 -421 233
rect -479 -183 -467 183
rect -433 -183 -421 183
rect 421 183 479 233
rect -479 -233 -421 -183
rect 421 -183 433 183
rect 467 -183 479 183
rect 421 -233 479 -183
rect -479 -245 479 -233
rect -479 -279 -371 -245
rect 371 -279 479 -245
rect -479 -291 479 -279
<< mvpsubdiffcont >>
rect -371 245 371 279
rect -467 -183 -433 183
rect 433 -183 467 183
rect -371 -279 371 -245
<< poly >>
rect -287 141 -187 157
rect -287 107 -271 141
rect -203 107 -187 141
rect -287 69 -187 107
rect -129 141 -29 157
rect -129 107 -113 141
rect -45 107 -29 141
rect -129 69 -29 107
rect 29 141 129 157
rect 29 107 45 141
rect 113 107 129 141
rect 29 69 129 107
rect 187 141 287 157
rect 187 107 203 141
rect 271 107 287 141
rect 187 69 287 107
rect -287 -157 -187 -131
rect -129 -157 -29 -131
rect 29 -157 129 -131
rect 187 -157 287 -131
<< polycont >>
rect -271 107 -203 141
rect -113 107 -45 141
rect 45 107 113 141
rect 203 107 271 141
<< locali >>
rect -467 245 -371 279
rect 371 245 467 279
rect -467 183 -433 245
rect 433 183 467 245
rect -287 107 -271 141
rect -203 107 -187 141
rect -129 107 -113 141
rect -45 107 -29 141
rect 29 107 45 141
rect 113 107 129 141
rect 187 107 203 141
rect 271 107 287 141
rect -333 57 -299 73
rect -333 -135 -299 -119
rect -175 57 -141 73
rect -175 -135 -141 -119
rect -17 57 17 73
rect -17 -135 17 -119
rect 141 57 175 73
rect 141 -135 175 -119
rect 299 57 333 73
rect 299 -135 333 -119
rect -467 -279 -433 -183
rect 433 -279 467 -183
<< viali >>
rect -271 107 -203 141
rect -113 107 -45 141
rect 45 107 113 141
rect 203 107 271 141
rect -333 -102 -299 -32
rect -175 -30 -141 40
rect -17 -102 17 -32
rect 141 -30 175 40
rect 299 -102 333 -32
rect -433 -279 -371 -245
rect -371 -279 371 -245
rect 371 -279 433 -245
<< metal1 >>
rect -283 141 -191 147
rect -283 107 -271 141
rect -203 107 -191 141
rect -283 101 -191 107
rect -125 141 -33 147
rect -125 107 -113 141
rect -45 107 -33 141
rect -125 101 -33 107
rect 33 141 125 147
rect 33 107 45 141
rect 113 107 125 141
rect 33 101 125 107
rect 191 141 283 147
rect 191 107 203 141
rect 271 107 283 141
rect 191 101 283 107
rect -181 40 -135 52
rect -339 -32 -293 -20
rect -339 -102 -333 -32
rect -299 -102 -293 -32
rect -181 -30 -175 40
rect -141 -30 -135 40
rect 135 40 181 52
rect -181 -42 -135 -30
rect -23 -32 23 -20
rect -339 -114 -293 -102
rect -23 -102 -17 -32
rect 17 -102 23 -32
rect 135 -30 141 40
rect 175 -30 181 40
rect 135 -42 181 -30
rect 293 -32 339 -20
rect -23 -114 23 -102
rect 293 -102 299 -32
rect 333 -102 339 -32
rect 293 -114 339 -102
rect -445 -245 445 -239
rect -445 -279 -433 -245
rect 433 -279 445 -245
rect -445 -285 445 -279
<< properties >>
string FIXED_BBOX -450 -262 450 262
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.50 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -40 viadrn +40 viagate 100 viagb 100 viagr 0 viagl 0 viagt 0
<< end >>
