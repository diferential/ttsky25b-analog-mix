magic
tech sky130A
magscale 1 2
timestamp 1762741441
<< pwell >>
rect -325 -1213 325 1213
<< nmoslvt >>
rect -129 603 -29 1003
rect 29 603 129 1003
rect -129 47 -29 447
rect 29 47 129 447
rect -129 -509 -29 -109
rect 29 -509 129 -109
rect -129 -1065 -29 -665
rect 29 -1065 129 -665
<< ndiff >>
rect -187 991 -129 1003
rect -187 615 -175 991
rect -141 615 -129 991
rect -187 603 -129 615
rect -29 991 29 1003
rect -29 615 -17 991
rect 17 615 29 991
rect -29 603 29 615
rect 129 991 187 1003
rect 129 615 141 991
rect 175 615 187 991
rect 129 603 187 615
rect -187 435 -129 447
rect -187 59 -175 435
rect -141 59 -129 435
rect -187 47 -129 59
rect -29 435 29 447
rect -29 59 -17 435
rect 17 59 29 435
rect -29 47 29 59
rect 129 435 187 447
rect 129 59 141 435
rect 175 59 187 435
rect 129 47 187 59
rect -187 -121 -129 -109
rect -187 -497 -175 -121
rect -141 -497 -129 -121
rect -187 -509 -129 -497
rect -29 -121 29 -109
rect -29 -497 -17 -121
rect 17 -497 29 -121
rect -29 -509 29 -497
rect 129 -121 187 -109
rect 129 -497 141 -121
rect 175 -497 187 -121
rect 129 -509 187 -497
rect -187 -677 -129 -665
rect -187 -1053 -175 -677
rect -141 -1053 -129 -677
rect -187 -1065 -129 -1053
rect -29 -677 29 -665
rect -29 -1053 -17 -677
rect 17 -1053 29 -677
rect -29 -1065 29 -1053
rect 129 -677 187 -665
rect 129 -1053 141 -677
rect 175 -1053 187 -677
rect 129 -1065 187 -1053
<< ndiffc >>
rect -175 615 -141 991
rect -17 615 17 991
rect 141 615 175 991
rect -175 59 -141 435
rect -17 59 17 435
rect 141 59 175 435
rect -175 -497 -141 -121
rect -17 -497 17 -121
rect 141 -497 175 -121
rect -175 -1053 -141 -677
rect -17 -1053 17 -677
rect 141 -1053 175 -677
<< psubdiff >>
rect -289 1143 -193 1177
rect 193 1143 289 1177
rect -289 1081 -255 1143
rect 255 1081 289 1143
rect -289 -1143 -255 -1081
rect 255 -1143 289 -1081
rect -289 -1177 -193 -1143
rect 193 -1177 289 -1143
<< psubdiffcont >>
rect -193 1143 193 1177
rect -289 -1081 -255 1081
rect 255 -1081 289 1081
rect -193 -1177 193 -1143
<< poly >>
rect -129 1075 -29 1091
rect -129 1041 -113 1075
rect -45 1041 -29 1075
rect -129 1003 -29 1041
rect 29 1075 129 1091
rect 29 1041 45 1075
rect 113 1041 129 1075
rect 29 1003 129 1041
rect -129 577 -29 603
rect 29 577 129 603
rect -129 519 -29 535
rect -129 485 -113 519
rect -45 485 -29 519
rect -129 447 -29 485
rect 29 519 129 535
rect 29 485 45 519
rect 113 485 129 519
rect 29 447 129 485
rect -129 21 -29 47
rect 29 21 129 47
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -109 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -109 129 -71
rect -129 -535 -29 -509
rect 29 -535 129 -509
rect -129 -593 -29 -577
rect -129 -627 -113 -593
rect -45 -627 -29 -593
rect -129 -665 -29 -627
rect 29 -593 129 -577
rect 29 -627 45 -593
rect 113 -627 129 -593
rect 29 -665 129 -627
rect -129 -1091 -29 -1065
rect 29 -1091 129 -1065
<< polycont >>
rect -113 1041 -45 1075
rect 45 1041 113 1075
rect -113 485 -45 519
rect 45 485 113 519
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect -113 -627 -45 -593
rect 45 -627 113 -593
<< locali >>
rect -289 1143 -193 1177
rect 193 1143 289 1177
rect -289 1081 -255 1143
rect 255 1081 289 1143
rect -129 1041 -113 1075
rect -45 1041 -29 1075
rect 29 1041 45 1075
rect 113 1041 129 1075
rect -175 991 -141 1007
rect -175 599 -141 615
rect -17 991 17 1007
rect -17 599 17 615
rect 141 991 175 1007
rect 141 599 175 615
rect -129 485 -113 519
rect -45 485 -29 519
rect 29 485 45 519
rect 113 485 129 519
rect -175 435 -141 451
rect -175 43 -141 59
rect -17 435 17 451
rect -17 43 17 59
rect 141 435 175 451
rect 141 43 175 59
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect -175 -121 -141 -105
rect -175 -513 -141 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 141 -121 175 -105
rect 141 -513 175 -497
rect -129 -627 -113 -593
rect -45 -627 -29 -593
rect 29 -627 45 -593
rect 113 -627 129 -593
rect -175 -677 -141 -661
rect -175 -1069 -141 -1053
rect -17 -677 17 -661
rect -17 -1069 17 -1053
rect 141 -677 175 -661
rect 141 -1069 175 -1053
rect -289 -1143 -255 -1081
rect 255 -1143 289 -1081
rect -289 -1177 -193 -1143
rect 193 -1177 289 -1143
<< viali >>
rect -102 1143 102 1177
rect -113 1041 -45 1075
rect 45 1041 113 1075
rect -175 632 -141 782
rect -17 824 17 974
rect 141 632 175 782
rect -113 485 -45 519
rect 45 485 113 519
rect -289 -457 -255 457
rect -175 76 -141 226
rect -17 268 17 418
rect 141 76 175 226
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect -175 -480 -141 -330
rect -17 -288 17 -138
rect 141 -480 175 -330
rect 255 -457 289 457
rect -113 -627 -45 -593
rect 45 -627 113 -593
rect -175 -1036 -141 -886
rect -17 -844 17 -694
rect 141 -1036 175 -886
rect -102 -1177 102 -1143
<< metal1 >>
rect -114 1177 114 1183
rect -114 1143 -102 1177
rect 102 1143 114 1177
rect -114 1137 114 1143
rect -125 1075 -33 1081
rect -125 1041 -113 1075
rect -45 1041 -33 1075
rect -125 1035 -33 1041
rect 33 1075 125 1081
rect 33 1041 45 1075
rect 113 1041 125 1075
rect 33 1035 125 1041
rect -23 974 23 986
rect -23 824 -17 974
rect 17 824 23 974
rect -23 812 23 824
rect -181 782 -135 794
rect -181 632 -175 782
rect -141 632 -135 782
rect -181 620 -135 632
rect 135 782 181 794
rect 135 632 141 782
rect 175 632 181 782
rect 135 620 181 632
rect -125 519 -33 525
rect -125 485 -113 519
rect -45 485 -33 519
rect -125 479 -33 485
rect 33 519 125 525
rect 33 485 45 519
rect 113 485 125 519
rect 33 479 125 485
rect -295 457 -249 469
rect -295 -457 -289 457
rect -255 -457 -249 457
rect 249 457 295 469
rect -23 418 23 430
rect -23 268 -17 418
rect 17 268 23 418
rect -23 256 23 268
rect -181 226 -135 238
rect -181 76 -175 226
rect -141 76 -135 226
rect -181 64 -135 76
rect 135 226 181 238
rect 135 76 141 226
rect 175 76 181 226
rect 135 64 181 76
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect -23 -138 23 -126
rect -23 -288 -17 -138
rect 17 -288 23 -138
rect -23 -300 23 -288
rect -295 -469 -249 -457
rect -181 -330 -135 -318
rect -181 -480 -175 -330
rect -141 -480 -135 -330
rect -181 -492 -135 -480
rect 135 -330 181 -318
rect 135 -480 141 -330
rect 175 -480 181 -330
rect 249 -457 255 457
rect 289 -457 295 457
rect 249 -469 295 -457
rect 135 -492 181 -480
rect -125 -593 -33 -587
rect -125 -627 -113 -593
rect -45 -627 -33 -593
rect -125 -633 -33 -627
rect 33 -593 125 -587
rect 33 -627 45 -593
rect 113 -627 125 -593
rect 33 -633 125 -627
rect -23 -694 23 -682
rect -23 -844 -17 -694
rect 17 -844 23 -694
rect -23 -856 23 -844
rect -181 -886 -135 -874
rect -181 -1036 -175 -886
rect -141 -1036 -135 -886
rect -181 -1048 -135 -1036
rect 135 -886 181 -874
rect 135 -1036 141 -886
rect 175 -1036 181 -886
rect 135 -1048 181 -1036
rect -114 -1143 114 -1137
rect -114 -1177 -102 -1143
rect 102 -1177 114 -1143
rect -114 -1183 114 -1177
<< properties >>
string FIXED_BBOX -272 -1160 272 1160
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.5 m 4 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -40 viadrn +40 viagate 100 viagb 40 viagr 40 viagl 40 viagt 40
string sky130_fd_pr__nfet_01v8_lvt_GXPBWL parameters
<< end >>
