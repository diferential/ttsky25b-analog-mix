magic
tech sky130A
magscale 1 2
timestamp 1725635217
<< pwell >>
rect -515 -658 515 658
<< mvnmos >>
rect -287 -400 -187 400
rect -129 -400 -29 400
rect 29 -400 129 400
rect 187 -400 287 400
<< mvndiff >>
rect -345 388 -287 400
rect -345 -388 -333 388
rect -299 -388 -287 388
rect -345 -400 -287 -388
rect -187 388 -129 400
rect -187 -388 -175 388
rect -141 -388 -129 388
rect -187 -400 -129 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 129 388 187 400
rect 129 -388 141 388
rect 175 -388 187 388
rect 129 -400 187 -388
rect 287 388 345 400
rect 287 -388 299 388
rect 333 -388 345 388
rect 287 -400 345 -388
<< mvndiffc >>
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
<< mvpsubdiff >>
rect -479 610 479 622
rect -479 576 -371 610
rect 371 576 479 610
rect -479 564 479 576
rect -479 514 -421 564
rect -479 -514 -467 514
rect -433 -514 -421 514
rect 421 514 479 564
rect -479 -564 -421 -514
rect 421 -514 433 514
rect 467 -514 479 514
rect 421 -564 479 -514
rect -479 -576 479 -564
rect -479 -610 -371 -576
rect 371 -610 479 -576
rect -479 -622 479 -610
<< mvpsubdiffcont >>
rect -371 576 371 610
rect -467 -514 -433 514
rect 433 -514 467 514
rect -371 -610 371 -576
<< poly >>
rect -287 472 -187 488
rect -287 438 -271 472
rect -203 438 -187 472
rect -287 400 -187 438
rect -129 472 -29 488
rect -129 438 -113 472
rect -45 438 -29 472
rect -129 400 -29 438
rect 29 472 129 488
rect 29 438 45 472
rect 113 438 129 472
rect 29 400 129 438
rect 187 472 287 488
rect 187 438 203 472
rect 271 438 287 472
rect 187 400 287 438
rect -287 -438 -187 -400
rect -287 -472 -271 -438
rect -203 -472 -187 -438
rect -287 -488 -187 -472
rect -129 -438 -29 -400
rect -129 -472 -113 -438
rect -45 -472 -29 -438
rect -129 -488 -29 -472
rect 29 -438 129 -400
rect 29 -472 45 -438
rect 113 -472 129 -438
rect 29 -488 129 -472
rect 187 -438 287 -400
rect 187 -472 203 -438
rect 271 -472 287 -438
rect 187 -488 287 -472
<< polycont >>
rect -271 438 -203 472
rect -113 438 -45 472
rect 45 438 113 472
rect 203 438 271 472
rect -271 -472 -203 -438
rect -113 -472 -45 -438
rect 45 -472 113 -438
rect 203 -472 271 -438
<< locali >>
rect -467 576 -371 610
rect 371 576 467 610
rect -467 514 -433 576
rect 433 514 467 576
rect -287 438 -271 472
rect -203 438 -187 472
rect -129 438 -113 472
rect -45 438 -29 472
rect 29 438 45 472
rect 113 438 129 472
rect 187 438 203 472
rect 271 438 287 472
rect -333 388 -299 404
rect -333 -404 -299 -388
rect -175 388 -141 404
rect -175 -404 -141 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 141 388 175 404
rect 141 -404 175 -388
rect 299 388 333 404
rect 299 -404 333 -388
rect -287 -472 -271 -438
rect -203 -472 -187 -438
rect -129 -472 -113 -438
rect -45 -472 -29 -438
rect 29 -472 45 -438
rect 113 -472 129 -438
rect 187 -472 203 -438
rect 271 -472 287 -438
rect -467 -576 -433 -514
rect 433 -576 467 -514
rect -467 -610 -371 -576
rect 371 -610 467 -576
<< viali >>
rect -271 438 -203 472
rect -113 438 -45 472
rect 45 438 113 472
rect 203 438 271 472
rect -467 -230 -433 230
rect -333 -155 -299 155
rect -175 61 -141 371
rect -17 -155 17 155
rect 141 61 175 371
rect 299 -155 333 155
rect 433 -230 467 230
rect -271 -472 -203 -438
rect -113 -472 -45 -438
rect 45 -472 113 -438
rect 203 -472 271 -438
rect -173 -610 173 -576
<< metal1 >>
rect -283 472 -191 478
rect -283 438 -271 472
rect -203 438 -191 472
rect -283 432 -191 438
rect -125 472 -33 478
rect -125 438 -113 472
rect -45 438 -33 472
rect -125 432 -33 438
rect 33 472 125 478
rect 33 438 45 472
rect 113 438 125 472
rect 33 432 125 438
rect 191 472 283 478
rect 191 438 203 472
rect 271 438 283 472
rect 191 432 283 438
rect -181 371 -135 383
rect -473 230 -427 242
rect -473 -230 -467 230
rect -433 -230 -427 230
rect -339 155 -293 167
rect -339 -155 -333 155
rect -299 -155 -293 155
rect -181 61 -175 371
rect -141 61 -135 371
rect 135 371 181 383
rect -181 49 -135 61
rect -23 155 23 167
rect -339 -167 -293 -155
rect -23 -155 -17 155
rect 17 -155 23 155
rect 135 61 141 371
rect 175 61 181 371
rect 427 230 473 242
rect 135 49 181 61
rect 293 155 339 167
rect -23 -167 23 -155
rect 293 -155 299 155
rect 333 -155 339 155
rect 293 -167 339 -155
rect -473 -242 -427 -230
rect 427 -230 433 230
rect 467 -230 473 230
rect 427 -242 473 -230
rect -283 -438 -191 -432
rect -283 -472 -271 -438
rect -203 -472 -191 -438
rect -283 -478 -191 -472
rect -125 -438 -33 -432
rect -125 -472 -113 -438
rect -45 -472 -33 -438
rect -125 -478 -33 -472
rect 33 -438 125 -432
rect 33 -472 45 -438
rect 113 -472 125 -438
rect 33 -478 125 -472
rect 191 -438 283 -432
rect 191 -472 203 -438
rect 271 -472 283 -438
rect 191 -478 283 -472
rect -185 -576 185 -570
rect -185 -610 -173 -576
rect 173 -610 185 -576
rect -185 -616 185 -610
<< properties >>
string FIXED_BBOX -450 -593 450 593
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -40 viadrn 40 viagate 100 viagb 40 viagr 40 viagl 40 viagt 0
string sky130_fd_pr__nfet_g5v0d10v5_R4FM4P parameters
<< end >>
