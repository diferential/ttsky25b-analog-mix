magic
tech sky130A
magscale 1 2
timestamp 1762742125
<< viali >>
rect 860 2600 1360 2660
rect 860 2360 1360 2420
rect 720 1720 1220 1780
<< metal1 >>
rect 2440 3500 4920 3620
rect 2440 3420 3680 3500
rect 160 2760 600 3160
rect 1910 3000 1920 3140
rect 2060 3000 2070 3140
rect 1910 2760 1920 2900
rect 2060 2760 2070 2900
rect 2440 2860 2620 3420
rect 3940 3380 4560 3440
rect 2700 3020 2760 3040
rect 3000 3020 3060 3120
rect 3110 3100 3120 3180
rect 3500 3100 3510 3180
rect 3780 3020 3860 3026
rect 2690 2940 2700 3020
rect 2780 2940 2790 3020
rect 2970 2940 2980 3020
rect 3060 2940 3070 3020
rect 3310 2940 3320 3020
rect 3500 2940 3510 3020
rect 2440 2780 2460 2860
rect 2580 2780 2620 2860
rect 848 2660 1372 2666
rect 80 2600 860 2660
rect 1360 2600 2000 2660
rect 80 2420 2000 2600
rect 2440 2480 2620 2780
rect 80 2360 860 2420
rect 1360 2360 2000 2420
rect 848 2354 1372 2360
rect 2280 2280 2620 2480
rect 200 1880 640 2280
rect 1550 2120 1560 2260
rect 1700 2120 1710 2260
rect 1550 1880 1560 2020
rect 1700 1880 1710 2020
rect 730 1786 740 1800
rect 708 1780 740 1786
rect 940 1786 950 1800
rect 940 1780 1232 1786
rect 708 1720 720 1780
rect 1220 1720 1232 1780
rect 708 1714 1232 1720
rect 0 1520 660 1540
rect 0 1420 340 1520
rect 480 1420 660 1520
rect 0 1240 660 1420
rect 2280 1360 2480 2280
rect 2700 2040 2760 2940
rect 3000 2840 3060 2940
rect 3110 2780 3120 2860
rect 3500 2780 3510 2860
rect 2630 1960 2640 2040
rect 2740 1960 2760 2040
rect 3040 2340 3700 2440
rect 3040 1680 3120 2340
rect 3180 2220 3540 2260
rect 3170 2160 3180 2220
rect 3240 2160 3480 2220
rect 3540 2160 3550 2220
rect 3180 2140 3540 2160
rect 3310 1920 3320 2060
rect 3420 1920 3430 2060
rect 3230 1780 3240 1840
rect 3500 1780 3510 1840
rect 3620 1680 3700 2340
rect 3780 2040 3860 2940
rect 3940 2540 4020 3380
rect 4370 3160 4380 3260
rect 4480 3160 4490 3260
rect 4700 3060 4920 3500
rect 4240 2940 4920 3060
rect 4700 2840 4920 2940
rect 4120 2620 4920 2840
rect 3940 2480 4560 2540
rect 3770 1960 3780 2040
rect 3860 1960 3870 2040
rect 3040 1560 3740 1680
rect 3040 1160 3120 1560
rect 3320 1280 3420 1500
rect 3230 1220 3240 1280
rect 3500 1220 3510 1280
rect 3620 1160 3740 1560
rect 3040 1040 3740 1160
rect 0 560 80 640
rect 3040 600 3120 1040
rect 3320 720 3420 940
rect 3230 660 3240 720
rect 3500 660 3510 720
rect 3620 600 3740 1040
rect 3940 1660 4020 2480
rect 4370 2240 4380 2340
rect 4480 2240 4490 2340
rect 4700 2160 4920 2620
rect 4240 2040 4920 2160
rect 4700 1960 4920 2040
rect 4120 1740 4920 1960
rect 3940 1600 4560 1660
rect 3940 770 4020 1600
rect 4370 1380 4380 1480
rect 4480 1380 4490 1480
rect 4700 1300 4920 1740
rect 4240 1180 4920 1300
rect 4700 1060 4920 1180
rect 4120 840 4920 1060
rect 3930 700 3940 770
rect 4020 760 4030 770
rect 4020 700 4560 760
rect 2680 480 3740 600
rect 4380 560 4460 700
rect 770 80 780 100
rect 20 0 780 80
rect 880 80 890 100
rect 2680 80 3120 480
rect 3310 240 3320 380
rect 3420 240 3430 380
rect 3230 120 3240 180
rect 3500 120 3510 180
rect 3620 80 3740 480
rect 4700 420 4920 840
rect 880 0 3740 80
rect 20 -40 3740 0
rect 4040 -40 4920 420
<< via1 >>
rect 1920 3000 2060 3140
rect 1920 2760 2060 2900
rect 3120 3100 3500 3180
rect 2700 2940 2780 3020
rect 2980 2940 3060 3020
rect 3320 2940 3500 3020
rect 3780 2940 3860 3020
rect 2460 2780 2580 2860
rect 1560 2120 1700 2260
rect 1560 1880 1700 2020
rect 740 1780 940 1800
rect 740 1720 940 1780
rect 340 1420 480 1520
rect 3120 2780 3500 2860
rect 2640 1960 2740 2040
rect 3180 2160 3240 2220
rect 3480 2160 3540 2220
rect 3320 1920 3420 2060
rect 3240 1780 3500 1840
rect 4380 3160 4480 3260
rect 3780 1960 3860 2040
rect 3240 1220 3500 1280
rect 3240 660 3500 720
rect 4380 2240 4480 2340
rect 4380 1380 4480 1480
rect 3940 700 4020 770
rect 780 0 880 100
rect 3320 240 3420 380
rect 3240 120 3500 180
<< metal2 >>
rect 4380 3260 4480 3270
rect 3120 3180 3500 3190
rect 1900 3140 3120 3180
rect 1900 3000 1920 3140
rect 2060 3100 3120 3140
rect 4380 3150 4480 3160
rect 2060 3000 2080 3100
rect 3120 3090 3500 3100
rect 1900 2980 2080 3000
rect 2700 3020 2780 3030
rect 2940 3020 3060 3030
rect 2780 2940 2980 3020
rect 2700 2930 2780 2940
rect 2940 2930 3060 2940
rect 1900 2900 2080 2920
rect 2940 2910 3040 2930
rect 1900 2760 1920 2900
rect 2060 2860 2620 2900
rect 2060 2780 2460 2860
rect 2580 2780 2620 2860
rect 2060 2760 2620 2780
rect 3120 2870 3200 3090
rect 3320 3020 3500 3030
rect 3500 2940 3780 3020
rect 3860 2940 3866 3020
rect 3320 2930 3500 2940
rect 3120 2860 3500 2870
rect 3120 2770 3500 2780
rect 1900 2740 2620 2760
rect 4380 2340 4480 2350
rect 1560 2260 1700 2270
rect 1700 2220 3560 2260
rect 4380 2230 4480 2240
rect 1700 2160 3180 2220
rect 3240 2160 3480 2220
rect 3540 2160 3560 2220
rect 1700 2140 3560 2160
rect 1560 2110 1700 2120
rect 3320 2060 3420 2070
rect 2640 2040 2740 2050
rect 1560 2020 1700 2030
rect 340 1880 1560 2000
rect 340 1520 480 1880
rect 1560 1870 1700 1880
rect 340 1410 480 1420
rect 740 1800 940 1810
rect 740 100 940 1720
rect 2640 810 2740 1960
rect 2960 1960 3320 2040
rect 2960 1280 3040 1960
rect 3780 2040 3860 2050
rect 3420 1960 3780 2040
rect 3780 1950 3860 1960
rect 3320 1910 3420 1920
rect 3240 1840 3500 1850
rect 3500 1780 3900 1840
rect 3240 1770 3500 1780
rect 4380 1480 4480 1490
rect 4380 1370 4480 1380
rect 3240 1280 3500 1290
rect 2960 1220 3240 1280
rect 2960 720 3040 1220
rect 3240 1210 3500 1220
rect 3940 770 4020 780
rect 3240 720 3500 730
rect 2960 660 3240 720
rect 2960 180 3040 660
rect 3240 650 3500 660
rect 3940 420 4020 700
rect 3320 380 4020 420
rect 3420 340 4020 380
rect 3320 230 3420 240
rect 3240 180 3500 190
rect 2960 120 3240 180
rect 3240 110 3500 120
rect 740 0 780 100
rect 880 0 940 100
rect 740 -40 940 0
use lvl_shift_lohi1  lvl_shift_lohi1_0
timestamp 1762742125
transform 1 0 0 0 1 0
box 0 0 2820 1680
use sky130_fd_pr__nfet_01v8_lvt_GXPBWL  sky130_fd_pr__nfet_01v8_lvt_GXPBWL_0
timestamp 1762742125
transform -1 0 3365 0 -1 1213
box -325 -1213 325 1213
use sky130_fd_pr__nfet_g5v0d10v5_FLD2WH  sky130_fd_pr__nfet_g5v0d10v5_FLD2WH_0
timestamp 1762742125
transform 0 -1 3267 1 0 2977
box -357 -427 357 427
use sky130_fd_pr__pfet_g5v0d10v5_PY9F4X  sky130_fd_pr__pfet_g5v0d10v5_PY9F4X_0
timestamp 1762742125
transform 1 0 4427 0 1 2262
box -387 -462 387 462
use sky130_fd_pr__pfet_g5v0d10v5_PY9F4X  sky130_fd_pr__pfet_g5v0d10v5_PY9F4X_1
timestamp 1762742125
transform 1 0 4427 0 1 482
box -387 -462 387 462
use sky130_fd_pr__pfet_g5v0d10v5_PY9F4X  sky130_fd_pr__pfet_g5v0d10v5_PY9F4X_2
timestamp 1762742125
transform 1 0 4427 0 1 1382
box -387 -462 387 462
use sky130_fd_pr__pfet_g5v0d10v5_PY9F4X  sky130_fd_pr__pfet_g5v0d10v5_PY9F4X_3
timestamp 1762742125
transform 1 0 4427 0 1 3162
box -387 -462 387 462
use sky130_fd_pr__res_high_po_0p69_SYH6D8  sky130_fd_pr__res_high_po_0p69_SYH6D8_0
timestamp 1762742125
transform 0 1 1038 -1 0 2072
box -352 -998 352 998
use sky130_fd_pr__res_xhigh_po_0p69_A2KNKC  sky130_fd_pr__res_xhigh_po_0p69_A2KNKC_0
timestamp 1762742125
transform 0 -1 1198 1 0 2952
box -352 -1198 352 1198
<< labels >>
flabel metal1 0 560 80 640 0 FreeSans 800 0 0 0 EN_RESH
port 0 nsew
flabel metal2 3840 1780 3900 1840 0 FreeSans 800 0 0 0 EN_RESL
port 1 nsew
flabel metal2 4380 3160 4480 3260 0 FreeSans 800 0 0 0 VOUT1
port 2 nsew
flabel metal2 4380 2240 4480 2340 0 FreeSans 800 0 0 0 VOUT2
port 3 nsew
flabel metal2 4380 1380 4480 1480 0 FreeSans 800 0 0 0 VOUT3
port 4 nsew
flabel metal1 2440 3420 2640 3620 0 FreeSans 800 0 0 0 VDDH
port 5 nsew
flabel metal1 0 1340 200 1540 0 FreeSans 800 0 0 0 VDDL
port 6 nsew
flabel metal1 2720 -40 2880 120 0 FreeSans 800 0 0 0 VSS
port 7 nsew
flabel metal2 2960 1960 3040 2040 0 FreeSans 800 0 0 0 VMID
<< end >>
