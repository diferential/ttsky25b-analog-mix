magic
tech sky130A
magscale 1 2
timestamp 1762800570
<< pwell >>
rect 16800 2270 18200 3080
rect 16800 2260 17180 2270
rect 17270 2260 18200 2270
rect 16800 1920 18200 2260
<< mvpsubdiff >>
rect 17320 3000 17760 3040
rect 16840 2920 17360 3000
rect 17720 2920 18160 3000
rect 16840 2040 16920 2920
rect 17320 2880 17760 2920
rect 18080 2040 18160 2920
rect 16840 1960 18160 2040
<< mvpsubdiffcont >>
rect 17360 2920 17720 3000
<< poly >>
rect 17170 2720 17260 2730
rect 17170 2670 17190 2720
rect 17240 2670 17260 2720
rect 17170 2650 17260 2670
rect 17550 2720 17640 2730
rect 17550 2670 17570 2720
rect 17620 2670 17640 2720
rect 17550 2650 17640 2670
rect 17200 2550 17230 2650
rect 17580 2580 17610 2650
rect 17310 2170 17340 2240
rect 17690 2170 17720 2240
rect 17280 2150 17370 2170
rect 17280 2100 17300 2150
rect 17350 2100 17370 2150
rect 17280 2090 17370 2100
rect 17660 2150 17750 2170
rect 17660 2100 17680 2150
rect 17730 2100 17750 2150
rect 17660 2090 17750 2100
<< polycont >>
rect 17190 2670 17240 2720
rect 17570 2670 17620 2720
rect 17300 2100 17350 2150
rect 17680 2100 17730 2150
<< locali >>
rect 17320 3000 17760 3040
rect 17320 2920 17360 3000
rect 17720 2920 17760 3000
rect 17320 2880 17760 2920
rect 17170 2720 17260 2730
rect 17170 2670 17190 2720
rect 17240 2670 17260 2720
rect 17170 2650 17260 2670
rect 17550 2720 17640 2730
rect 17550 2670 17570 2720
rect 17620 2670 17640 2720
rect 17550 2650 17640 2670
rect 17280 2150 17370 2170
rect 17280 2100 17300 2150
rect 17350 2100 17370 2150
rect 17280 2090 17370 2100
rect 17660 2150 17750 2170
rect 17660 2100 17680 2150
rect 17730 2100 17750 2150
rect 17660 2090 17750 2100
<< viali >>
rect 17360 2920 17720 3000
rect 17190 2670 17240 2710
rect 17570 2670 17620 2710
rect 17300 2110 17350 2150
rect 17680 2110 17730 2150
<< metal1 >>
rect 23090 11500 23100 11700
rect 23600 11500 23610 11700
rect 20590 9300 20600 9600
rect 20900 9300 20910 9600
rect 20440 8600 20450 8680
rect 20540 8600 20780 8680
rect 20590 7800 20600 8100
rect 21200 7800 21210 8100
rect 24680 8000 25560 8140
rect 25200 7540 25560 8000
rect 24600 7500 25560 7540
rect 21070 7080 21080 7400
rect 21400 7080 21410 7400
rect 25200 6800 25560 7500
rect 21030 4440 21380 4520
rect 21030 4240 21040 4440
rect 21360 4400 21380 4440
rect 21360 4240 21370 4400
rect 17348 3000 17732 3006
rect 17348 2920 17360 3000
rect 17720 2920 17732 3000
rect 17348 2914 17732 2920
rect 17170 2660 17180 2720
rect 17240 2716 17250 2720
rect 17240 2664 17252 2716
rect 17240 2660 17250 2664
rect 17550 2660 17560 2720
rect 17620 2716 17630 2720
rect 17620 2664 17632 2716
rect 17620 2660 17630 2664
rect 17880 2480 19500 2520
rect 17805 2450 19500 2480
rect 17880 2420 19500 2450
rect 19600 2420 19740 2520
rect 20210 2340 20220 2380
rect 17880 2320 20220 2340
rect 17810 2290 20220 2320
rect 17880 2240 20220 2290
rect 20210 2200 20220 2240
rect 20360 2340 20370 2380
rect 20360 2240 20410 2340
rect 20360 2200 20370 2240
rect 17290 2156 17300 2160
rect 17288 2104 17300 2156
rect 17290 2100 17300 2104
rect 17360 2100 17370 2160
rect 17670 2156 17680 2160
rect 17668 2104 17680 2156
rect 17670 2100 17680 2104
rect 17740 2100 17750 2160
<< via1 >>
rect 23100 11500 23600 11700
rect 20600 9300 20900 9600
rect 20450 8600 20540 8680
rect 20600 7800 21200 8100
rect 21080 7080 21400 7400
rect 21040 4240 21360 4440
rect 17360 2920 17720 3000
rect 17180 2710 17240 2720
rect 17180 2670 17190 2710
rect 17190 2670 17240 2710
rect 17180 2660 17240 2670
rect 17560 2710 17620 2720
rect 17560 2670 17570 2710
rect 17570 2670 17620 2710
rect 17560 2660 17620 2670
rect 19500 2420 19600 2520
rect 20220 2200 20360 2380
rect 17300 2150 17360 2160
rect 17300 2110 17350 2150
rect 17350 2110 17360 2150
rect 17300 2100 17360 2110
rect 17680 2150 17740 2160
rect 17680 2110 17730 2150
rect 17730 2110 17740 2150
rect 17680 2100 17740 2110
<< metal2 >>
rect 23100 11700 23600 11710
rect 23100 11490 23600 11500
rect 25020 11300 25120 11310
rect 25020 11190 25120 11200
rect 24400 9880 24560 9890
rect 24400 9710 24560 9720
rect 20600 9600 20900 9610
rect 20600 9290 20900 9300
rect 20440 8690 20540 8700
rect 20440 8580 20540 8590
rect 20600 8100 21200 8110
rect 20600 7790 21200 7800
rect 21080 7400 21400 7410
rect 21080 7070 21400 7080
rect 27320 6590 27560 6700
rect 23805 6320 27565 6590
rect 20560 5820 21040 5900
rect 20560 4520 20640 5820
rect 19440 4440 20640 4520
rect 20760 5660 21040 5740
rect 17360 3000 17720 3010
rect 17360 2910 17720 2920
rect 17160 2760 17270 2770
rect 17270 2640 17280 2760
rect 17160 2630 17270 2640
rect 17430 2520 17490 2910
rect 17560 2760 17670 2770
rect 17540 2640 17560 2760
rect 17560 2630 17670 2640
rect 19440 2520 19735 4440
rect 20760 3960 20840 5660
rect 24420 5532 24660 5934
rect 25520 5545 25720 5640
rect 25520 5455 25605 5545
rect 25695 5455 25720 5545
rect 25520 5420 25720 5455
rect 21030 4440 21380 4520
rect 21030 4400 21040 4440
rect 21360 4400 21380 4440
rect 21040 4230 21360 4240
rect 19440 2420 19500 2520
rect 19600 2420 19735 2520
rect 17240 2180 17350 2190
rect 17660 2180 17770 2190
rect 17350 2160 17360 2180
rect 17350 2060 17360 2100
rect 17770 2060 17780 2180
rect 17240 2050 17350 2060
rect 17660 2050 17770 2060
rect 19440 1782 19735 2420
rect 20140 3880 20840 3960
rect 20140 2380 20420 3880
rect 27320 2400 27560 6320
rect 20140 2200 20220 2380
rect 20360 2200 20420 2380
rect 20140 1855 20420 2200
rect 27120 2240 27640 2400
rect 27120 1945 27174 2240
rect 27469 1945 27640 2240
rect 27120 1920 27640 1945
rect 19436 1497 19445 1782
rect 19730 1497 19739 1782
rect 20136 1585 20145 1855
rect 20415 1585 20424 1855
rect 20140 1580 20420 1585
rect 19440 1492 19735 1497
<< via2 >>
rect 23100 11500 23600 11700
rect 25020 11200 25120 11300
rect 24400 9720 24560 9880
rect 20600 9300 20900 9600
rect 20440 8680 20540 8690
rect 20440 8600 20450 8680
rect 20450 8600 20540 8680
rect 20440 8590 20540 8600
rect 20600 7800 21200 8100
rect 21080 7080 21400 7400
rect 17360 2920 17720 3000
rect 17160 2720 17270 2760
rect 17160 2660 17180 2720
rect 17180 2660 17240 2720
rect 17240 2660 17270 2720
rect 17160 2640 17270 2660
rect 17560 2720 17670 2760
rect 17560 2660 17620 2720
rect 17620 2660 17670 2720
rect 17560 2640 17670 2660
rect 25605 5455 25695 5545
rect 21040 4240 21360 4400
rect 17240 2160 17350 2180
rect 17240 2100 17300 2160
rect 17300 2100 17350 2160
rect 17240 2060 17350 2100
rect 17660 2160 17770 2180
rect 17660 2100 17680 2160
rect 17680 2100 17740 2160
rect 17740 2100 17770 2160
rect 17660 2060 17770 2100
rect 27174 1945 27469 2240
rect 19445 1497 19730 1782
rect 20145 1585 20415 1855
<< metal3 >>
rect 21640 41900 21960 42000
rect 13660 41899 21960 41900
rect 13660 41880 21681 41899
rect 13660 41700 13800 41880
rect 13790 41680 13800 41700
rect 13960 41701 21681 41880
rect 21879 41701 21960 41899
rect 13960 41700 21960 41701
rect 13960 41680 13970 41700
rect 21640 41640 21960 41700
rect 14470 41420 14480 41440
rect 14380 41240 14480 41420
rect 14640 41420 14650 41440
rect 22160 41420 22480 41520
rect 14640 41419 22480 41420
rect 14640 41240 22201 41419
rect 14380 41221 22201 41240
rect 22399 41221 22480 41419
rect 14380 41220 22480 41221
rect 22160 41160 22480 41220
rect 15110 41020 15120 41040
rect 14980 40840 15120 41020
rect 15280 41020 15290 41040
rect 22680 41020 23000 41120
rect 15280 41019 23000 41020
rect 15280 40840 22761 41019
rect 14980 40821 22761 40840
rect 22959 40821 23000 41019
rect 14980 40820 23000 40821
rect 22680 40760 23000 40820
rect 23200 40625 23520 40680
rect 15695 40624 23520 40625
rect 15695 40600 23281 40624
rect 15695 40415 15760 40600
rect 15750 40400 15760 40415
rect 15920 40416 23281 40600
rect 23489 40416 23520 40624
rect 15920 40415 23520 40416
rect 15920 40400 15930 40415
rect 23200 40320 23520 40415
rect 192 21586 198 21986
rect 598 21586 3360 21986
rect 794 20634 800 21034
rect 1200 20634 3360 21034
rect 20242 12118 20398 12122
rect 20242 12117 24098 12118
rect 20242 12116 23883 12117
rect 20398 11963 23883 12116
rect 24037 11963 24098 12117
rect 20398 11962 24098 11963
rect 20242 11956 20398 11962
rect 22600 11720 23800 11800
rect 22600 11420 22650 11720
rect 22960 11700 23800 11720
rect 22960 11500 23100 11700
rect 23600 11500 23800 11700
rect 22960 11420 23800 11500
rect 22600 11400 23800 11420
rect 25010 11300 25130 11305
rect 25580 11300 25720 11320
rect 25010 11200 25020 11300
rect 25120 11200 25600 11300
rect 25700 11200 25720 11300
rect 25010 11195 25130 11200
rect 25580 11180 25720 11200
rect 24390 9880 24570 9885
rect 24390 9720 24400 9880
rect 24560 9720 24570 9880
rect 24390 9715 24570 9720
rect 20590 9600 20910 9605
rect 244 9300 250 9600
rect 548 9300 20600 9600
rect 20900 9300 21200 9600
rect 20590 9295 20910 9300
rect 20242 8717 20838 8718
rect 20237 8563 20243 8717
rect 20397 8690 20838 8717
rect 20397 8590 20440 8690
rect 20540 8590 20838 8690
rect 20397 8563 20838 8590
rect 20242 8562 20838 8563
rect 20590 8100 21210 8105
rect 840 7800 850 8100
rect 1150 7800 20600 8100
rect 21200 7800 21210 8100
rect 20590 7795 21210 7800
rect 1401 7560 1799 7565
rect 1400 7559 5200 7560
rect 1400 7161 1401 7559
rect 1799 7440 5200 7559
rect 1799 7400 22600 7440
rect 1799 7161 21080 7400
rect 1400 7160 21080 7161
rect 1401 7155 1799 7160
rect 5000 7080 21080 7160
rect 21400 7080 22600 7400
rect 5000 7040 22600 7080
rect 22990 7400 23000 7430
rect 22990 7040 23600 7400
rect 25520 5549 25720 5640
rect 25520 5451 25601 5549
rect 25699 5451 25720 5549
rect 25520 5420 25720 5451
rect 801 4520 1199 4525
rect 800 4519 19960 4520
rect 800 4121 801 4519
rect 1199 4400 19960 4519
rect 20920 4400 21440 4560
rect 1199 4240 21040 4400
rect 21360 4240 21440 4400
rect 1199 4121 21440 4240
rect 800 4120 21440 4121
rect 801 4115 1199 4120
rect 17320 3000 17760 4120
rect 19600 4000 21440 4120
rect 17320 2920 17360 3000
rect 17720 2920 17760 3000
rect 17320 2880 17760 2920
rect 17150 2760 17280 2765
rect 14380 2640 14480 2760
rect 14680 2640 17160 2760
rect 17270 2640 17280 2760
rect 17150 2635 17280 2640
rect 17550 2760 17680 2765
rect 17550 2640 17560 2760
rect 17670 2640 17680 2760
rect 17550 2635 17680 2640
rect 17560 2440 17680 2635
rect 13740 2320 13800 2440
rect 14000 2320 17680 2440
rect 27169 2240 27474 2245
rect 17230 2180 17360 2185
rect 17230 2160 17240 2180
rect 15040 2040 15080 2160
rect 15280 2060 17240 2160
rect 17350 2060 17360 2180
rect 15280 2040 17360 2060
rect 17650 2180 17780 2185
rect 17650 2060 17660 2180
rect 17770 2060 17780 2180
rect 17650 2055 17780 2060
rect 17660 1760 17780 2055
rect 27169 1945 27174 2240
rect 27469 1945 27474 2240
rect 27169 1940 27474 1945
rect 20141 1860 20419 1865
rect 20140 1859 20420 1860
rect 19440 1786 19735 1787
rect 15680 1640 15760 1760
rect 15920 1640 17900 1760
rect 19435 1493 19441 1786
rect 19734 1493 19740 1786
rect 20140 1581 20141 1859
rect 20419 1581 20420 1859
rect 20140 1580 20420 1581
rect 27174 1744 27469 1940
rect 20141 1575 20419 1580
rect 19440 1492 19735 1493
rect 27174 1443 27469 1449
<< via3 >>
rect 13800 41680 13960 41880
rect 21681 41701 21879 41899
rect 14480 41240 14640 41440
rect 22201 41221 22399 41419
rect 15120 40840 15280 41040
rect 22761 40821 22959 41019
rect 15760 40400 15920 40600
rect 23281 40416 23489 40624
rect 198 21586 598 21986
rect 800 20634 1200 21034
rect 20242 11962 20398 12116
rect 23883 11963 24037 12117
rect 22650 11420 22960 11720
rect 25600 11200 25700 11300
rect 24400 9720 24560 9880
rect 250 9300 548 9600
rect 20243 8563 20397 8717
rect 850 7800 1150 8100
rect 1401 7161 1799 7559
rect 22600 7040 22990 7430
rect 25601 5545 25699 5549
rect 25601 5455 25605 5545
rect 25605 5455 25695 5545
rect 25695 5455 25699 5545
rect 25601 5451 25699 5455
rect 801 4121 1199 4519
rect 14480 2640 14680 2760
rect 13800 2320 14000 2440
rect 15080 2040 15280 2160
rect 15760 1640 15920 1760
rect 19441 1782 19734 1786
rect 19441 1497 19445 1782
rect 19445 1497 19730 1782
rect 19730 1497 19734 1782
rect 19441 1493 19734 1497
rect 20141 1855 20419 1859
rect 20141 1585 20145 1855
rect 20145 1585 20415 1855
rect 20415 1585 20419 1855
rect 20141 1581 20419 1585
rect 27174 1449 27469 1744
<< metal4 >>
rect 3006 44792 3066 45152
rect 3558 44792 3618 45152
rect 4110 44792 4170 45152
rect 4662 44792 4722 45152
rect 5214 44792 5274 45152
rect 5766 44792 5826 45152
rect 6318 44792 6378 45152
rect 6870 44792 6930 45152
rect 7422 44792 7482 45152
rect 7974 44792 8034 45152
rect 8526 44792 8586 45152
rect 9078 44792 9138 45152
rect 9630 44792 9690 45152
rect 10182 44792 10242 45152
rect 10734 44792 10794 45152
rect 11286 44792 11346 45152
rect 11838 44792 11898 45152
rect 12390 44792 12450 45152
rect 12942 44792 13002 45152
rect 13494 44792 13554 45152
rect 14046 44792 14106 45152
rect 14598 44792 14658 45152
rect 15150 44792 15210 45152
rect 15702 44792 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44840 19626 45152
rect 20118 44800 20178 45152
rect 20670 44800 20730 45152
rect 21222 44800 21282 45152
rect 960 44732 15762 44792
rect 960 44152 1020 44732
rect 6870 44722 6930 44732
rect 7974 44716 8034 44732
rect 15702 44730 15762 44732
rect 21774 44560 21834 45152
rect 22326 44560 22386 45152
rect 22878 44560 22938 45152
rect 23430 44560 23490 45152
rect 23982 44560 24042 45152
rect 24534 44560 24594 45152
rect 25086 44800 25146 45152
rect 25638 44800 25698 45152
rect 26190 44952 26250 45152
rect 200 21987 600 44152
rect 197 21986 600 21987
rect 197 21586 198 21986
rect 598 21586 600 21986
rect 197 21585 600 21586
rect 200 9600 600 21585
rect 800 21035 1200 44152
rect 799 21034 1201 21035
rect 799 20634 800 21034
rect 1200 20634 1201 21034
rect 799 20633 1201 20634
rect 200 9300 250 9600
rect 548 9300 600 9600
rect 200 1000 600 9300
rect 800 8100 1200 20633
rect 800 7800 850 8100
rect 1150 7800 1200 8100
rect 800 4519 1200 7800
rect 800 4121 801 4519
rect 1199 4121 1200 4519
rect 800 1000 1200 4121
rect 1400 20160 1800 44152
rect 13760 41880 14080 42560
rect 13760 41680 13800 41880
rect 13960 41680 14080 41880
rect 1400 19760 3360 20160
rect 1400 7559 1800 19760
rect 1400 7161 1401 7559
rect 1799 7161 1800 7559
rect 1400 1000 1800 7161
rect 13760 2440 14080 41680
rect 13760 2320 13800 2440
rect 14000 2320 14080 2440
rect 13760 2080 14080 2320
rect 14400 41440 14720 42560
rect 14400 41240 14480 41440
rect 14640 41240 14720 41440
rect 14400 2760 14720 41240
rect 15040 41040 15360 42560
rect 15040 41021 15120 41040
rect 15019 40840 15120 41021
rect 15280 40840 15360 41040
rect 15019 40819 15360 40840
rect 14400 2640 14480 2760
rect 14680 2640 14720 2760
rect 14400 2080 14720 2640
rect 15040 2160 15360 40819
rect 15040 2040 15080 2160
rect 15280 2040 15360 2160
rect 15040 1760 15360 2040
rect 15680 40600 16000 42560
rect 21680 42000 21880 44560
rect 21640 41899 21960 42000
rect 21640 41701 21681 41899
rect 21879 41701 21960 41899
rect 21640 41640 21960 41701
rect 15680 40400 15760 40600
rect 15920 40400 16000 40600
rect 21680 40420 21880 41640
rect 22200 41520 22400 44560
rect 22160 41419 22480 41520
rect 22160 41221 22201 41419
rect 22399 41221 22480 41419
rect 22160 41160 22480 41221
rect 22200 40420 22400 41160
rect 22760 41120 22960 44560
rect 22680 41019 23000 41120
rect 22680 40821 22761 41019
rect 22959 40821 23000 41019
rect 22680 40760 23000 40821
rect 22760 40420 22960 40760
rect 23280 40680 23490 44560
rect 23880 44410 24042 44560
rect 23880 43120 24040 44410
rect 24520 43280 24680 44560
rect 24400 43120 24680 43280
rect 23200 40624 23520 40680
rect 15680 1760 16000 40400
rect 23200 40416 23281 40624
rect 23489 40416 23520 40624
rect 23200 40320 23520 40416
rect 23882 12117 24038 43120
rect 20241 12116 20399 12117
rect 20241 11962 20242 12116
rect 20398 11962 20399 12116
rect 20241 11961 20399 11962
rect 23882 11963 23883 12117
rect 24037 11963 24038 12117
rect 20242 8717 20398 11961
rect 23882 11942 24038 11963
rect 20242 8563 20243 8717
rect 20397 8563 20398 8717
rect 20242 8562 20398 8563
rect 22600 11720 23000 11800
rect 22600 11420 22650 11720
rect 22960 11420 23000 11720
rect 22600 7431 23000 11420
rect 24400 9881 24560 43120
rect 25580 11300 25720 11320
rect 25580 11200 25600 11300
rect 25700 11200 25720 11300
rect 25580 11180 25720 11200
rect 24399 9880 24561 9881
rect 24399 9720 24400 9880
rect 24560 9720 24561 9880
rect 24399 9719 24561 9720
rect 22599 7430 23000 7431
rect 22599 7040 22600 7430
rect 22990 7040 23000 7430
rect 22599 7039 22991 7040
rect 25600 5640 25700 11180
rect 25520 5549 25720 5640
rect 25520 5451 25601 5549
rect 25699 5451 25720 5549
rect 25520 5420 25720 5451
rect 20140 1859 23600 1860
rect 15680 1640 15760 1760
rect 15920 1640 16000 1760
rect 15680 1600 16000 1640
rect 19440 1786 19735 1787
rect 19440 1493 19441 1786
rect 19734 1493 19735 1786
rect 20140 1581 20141 1859
rect 20419 1581 23600 1859
rect 20140 1580 23600 1581
rect 19440 440 19735 1493
rect 23320 440 23600 1580
rect 27173 1744 27470 1745
rect 27173 1449 27174 1744
rect 27469 1449 27470 1744
rect 27173 1448 27470 1449
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 440
rect 23370 0 23550 440
rect 27174 315 27469 1448
rect 27234 0 27414 315
use dram3t_charlie  dram3t_charlie_0
timestamp 1719885249
transform 1 0 17120 0 1 2240
box 0 0 720 340
use opamp3hvs  opamp3hvs_0
timestamp 1762794020
transform 1 0 20960 0 1 4240
box -1840 0 5400 3300
use root_currents1_3outs  root_currents1_3outs_0
timestamp 1762742125
transform 1 0 20640 0 1 8040
box 0 -40 4920 3624
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 1400 1000 1800 44152 1 FreeSans 1600 0 0 0 VAPWR
port 53 nsew power bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
