magic
tech sky130A
magscale 1 2
timestamp 1762740518
<< locali >>
rect -40 2900 4200 3020
rect -40 2880 2960 2900
rect -40 2540 100 2880
rect 1140 2720 2960 2880
rect 1140 2540 1280 2720
rect -40 2400 1280 2540
rect 120 2300 1280 2400
rect 2780 2560 2960 2720
rect 4000 2560 4200 2900
rect 2780 2280 4200 2560
rect -900 2180 -520 2240
rect -40 50 50 880
rect -40 40 4190 50
rect -40 20 4200 40
rect -40 -200 0 20
rect 60 -80 640 20
rect 700 -80 920 20
rect 980 -80 1200 20
rect 1260 -80 2580 20
rect 2640 -80 2860 20
rect 2920 -80 3140 20
rect 3200 -80 4080 20
rect 4140 -80 4200 20
rect 4160 -200 4200 -80
rect -40 -280 4200 -200
<< viali >>
rect 100 2540 1140 2880
rect 2960 2560 4000 2900
rect 0 -80 60 20
rect 640 -80 700 20
rect 920 -80 980 20
rect 1200 -80 1260 20
rect 2580 -80 2640 20
rect 2860 -80 2920 20
rect 3140 -80 3200 20
rect 4080 -80 4140 20
rect 0 -200 4160 -80
<< metal1 >>
rect -40 2960 4200 3020
rect -760 2760 -680 2920
rect -40 2900 2980 2960
rect 3080 2900 4200 2960
rect -40 2880 2960 2900
rect -40 2760 100 2880
rect -760 2680 100 2760
rect -900 2220 -860 2240
rect -980 2180 -800 2220
rect -980 2140 -820 2180
rect -980 1700 -860 2140
rect -760 2120 -680 2680
rect -40 2540 100 2680
rect 1140 2710 2960 2880
rect 1140 2540 1360 2710
rect 2680 2560 2960 2710
rect 4000 2560 4200 2900
rect 2680 2540 4200 2560
rect -40 2520 1390 2540
rect 2650 2520 4200 2540
rect -40 2400 4200 2520
rect 120 2300 4200 2400
rect 360 2280 440 2300
rect 730 2280 4200 2300
rect -800 1740 -640 2120
rect -980 1620 -820 1700
rect -600 1640 -560 2220
rect -980 1290 -900 1620
rect -500 1560 -420 2120
rect 1340 1810 1350 2070
rect 1410 1810 1420 2070
rect 1660 1810 1670 2070
rect 1730 1810 1740 2070
rect 1980 1810 1990 2070
rect 2050 1810 2060 2070
rect 2300 1810 2310 2070
rect 2370 1810 2380 2070
rect 2610 1810 2620 2070
rect 2680 1810 2690 2070
rect 4130 1880 4140 2040
rect 4320 1880 4330 2040
rect 840 1640 2680 1680
rect 160 1620 2680 1640
rect 160 1560 940 1620
rect -500 1520 940 1560
rect 1060 1600 2680 1620
rect 1060 1520 1120 1600
rect -500 1480 1120 1520
rect -500 1430 660 1480
rect -980 1210 230 1290
rect -40 400 50 880
rect 140 820 230 1210
rect 580 980 660 1430
rect 930 1260 990 1420
rect 1200 1340 1210 1420
rect 1270 1340 1280 1420
rect 920 1180 930 1260
rect 990 1180 1000 1260
rect 930 1050 990 1180
rect 1210 1050 1270 1340
rect 1480 1260 1540 1420
rect 1740 1340 1750 1420
rect 1810 1340 1820 1420
rect 2020 1340 2030 1420
rect 2090 1340 2100 1420
rect 1470 1180 1480 1260
rect 1540 1180 1550 1260
rect 1480 1050 1540 1180
rect 1750 1050 1810 1340
rect 2030 1050 2090 1340
rect 2310 1260 2370 1420
rect 2570 1340 2580 1420
rect 2640 1340 2650 1420
rect 2300 1180 2310 1260
rect 2370 1180 2380 1260
rect 2310 1050 2370 1180
rect 2580 1050 2640 1340
rect 2860 1260 2920 1420
rect 4140 1280 4320 1880
rect 2850 1180 2860 1260
rect 2920 1180 2930 1260
rect 2860 1050 2920 1180
rect 3420 1080 3460 1100
rect 570 900 580 980
rect 660 900 670 980
rect 130 740 140 820
rect 220 740 230 820
rect -40 80 160 400
rect 210 180 250 690
rect 280 590 350 610
rect 280 430 290 590
rect 280 420 350 430
rect 380 180 420 690
rect 190 120 200 180
rect 270 120 280 180
rect 350 120 360 180
rect 430 120 440 180
rect 380 110 420 120
rect 470 80 620 410
rect 830 280 840 440
rect 940 140 980 1050
rect 1110 900 1120 980
rect 1180 900 1190 980
rect 1010 740 1020 820
rect 1080 740 1090 820
rect 1220 140 1260 1050
rect 1490 140 1530 1050
rect 1650 900 1660 980
rect 1720 900 1730 980
rect 1560 740 1570 820
rect 1630 740 1640 820
rect 1760 140 1800 1050
rect 1830 280 1840 440
rect 2040 150 2080 1050
rect 2110 900 2120 980
rect 2180 900 2190 980
rect 2200 740 2210 820
rect 2270 740 2280 820
rect 2320 150 2360 1050
rect 2390 280 2400 440
rect 2590 150 2630 1050
rect 2670 900 2680 980
rect 2740 900 2750 980
rect 2760 740 2770 820
rect 2830 740 2840 820
rect 2870 150 2910 1050
rect 3410 1020 3460 1080
rect 3570 1080 3620 1100
rect 3080 640 3370 990
rect 3410 980 3450 1020
rect 3570 980 3610 1080
rect 3410 800 3440 980
rect 3470 830 3480 950
rect 3540 830 3550 950
rect 3580 800 3610 980
rect 3410 670 3450 800
rect 3570 680 3610 800
rect 3080 630 3320 640
rect 3080 550 3110 630
rect 3200 550 3320 630
rect 3380 550 3390 640
rect 3010 280 3020 440
rect 3080 220 3370 550
rect 3420 510 3460 670
rect -40 60 620 80
rect 3080 60 3340 220
rect 3410 180 3460 510
rect 3570 400 3600 680
rect 3630 440 3640 650
rect 3700 440 3710 650
rect 3570 180 3610 400
rect 3740 180 3780 1100
rect 3900 980 3940 1100
rect 4080 990 4320 1280
rect 3870 830 3880 950
rect 3910 800 3940 980
rect 3900 180 3940 800
rect 3990 640 4320 990
rect 3970 550 3980 640
rect 4040 550 4090 640
rect 4150 550 4320 640
rect 3990 220 4320 550
rect 3390 120 3400 180
rect 3470 120 3480 180
rect 3550 120 3560 180
rect 3630 120 3640 180
rect 3710 120 3720 180
rect 3790 120 3800 180
rect 3870 120 3880 180
rect 3950 120 3960 180
rect 4010 60 4320 220
rect -40 20 4320 60
rect -40 -200 0 20
rect 60 -80 640 20
rect 700 -80 920 20
rect 980 -80 1200 20
rect 1260 -80 2580 20
rect 2640 -80 2860 20
rect 2920 -80 3140 20
rect 3200 -80 4080 20
rect 4140 -80 4320 20
rect 4160 -200 4320 -80
rect -40 -280 4320 -200
<< via1 >>
rect 2980 2900 3080 2960
rect 2980 2740 3080 2900
rect 1350 1810 1410 2070
rect 1670 1810 1730 2070
rect 1990 1810 2050 2070
rect 2310 1810 2370 2070
rect 2620 1810 2680 2070
rect 4140 1880 4320 2040
rect 940 1520 1060 1620
rect 1210 1340 1270 1420
rect 930 1180 990 1260
rect 1750 1340 1810 1420
rect 2030 1340 2090 1420
rect 1480 1180 1540 1260
rect 2580 1340 2640 1420
rect 2310 1180 2370 1260
rect 2860 1180 2920 1260
rect 580 900 660 980
rect 140 740 220 820
rect 290 430 350 590
rect 200 120 270 180
rect 360 120 430 180
rect 840 280 900 440
rect 1120 900 1180 980
rect 1020 740 1080 820
rect 1300 280 1440 440
rect 1660 900 1720 980
rect 1570 740 1630 820
rect 1840 280 2000 440
rect 2120 900 2180 980
rect 2210 740 2270 820
rect 2400 280 2550 440
rect 2680 900 2740 980
rect 2770 740 2830 820
rect 3480 830 3540 950
rect 3110 550 3200 630
rect 3320 550 3380 640
rect 2950 280 3010 440
rect 3640 440 3700 650
rect 3810 830 3870 950
rect 3980 550 4040 640
rect 4090 550 4150 640
rect 3400 120 3470 180
rect 3560 120 3630 180
rect 3720 120 3790 180
rect 3880 120 3950 180
<< metal2 >>
rect 2980 2960 3080 2970
rect 2980 2730 3080 2740
rect 1350 2070 1410 2080
rect 1670 2070 1730 2080
rect 1990 2070 2050 2080
rect 2310 2070 2370 2080
rect 2620 2070 2680 2080
rect 1340 1810 1350 2070
rect 1410 1980 1670 2070
rect 1730 1980 1990 2070
rect 1410 1860 1660 1980
rect 1740 1860 1990 1980
rect 1410 1810 1670 1860
rect 1730 1810 1990 1860
rect 2050 1810 2310 2070
rect 2370 1810 2620 2070
rect 2680 1810 3660 2070
rect 4140 2040 4320 2050
rect 4140 1870 4320 1880
rect 1340 1800 3660 1810
rect 940 1620 1060 1630
rect 940 1510 1060 1520
rect 1210 1420 1270 1430
rect 1750 1420 1810 1430
rect 2030 1420 2090 1430
rect 2580 1420 2640 1430
rect -40 1340 1210 1420
rect 1270 1340 1750 1420
rect 1810 1340 2030 1420
rect 2090 1340 2580 1420
rect 2640 1340 3060 1420
rect 1210 1330 1270 1340
rect 1750 1330 1810 1340
rect 2030 1330 2090 1340
rect 2580 1330 2640 1340
rect 930 1260 990 1270
rect 1480 1260 1540 1270
rect 2310 1260 2370 1270
rect 2860 1260 2920 1270
rect -40 1180 930 1260
rect 990 1180 1480 1260
rect 1540 1180 2310 1260
rect 2370 1180 2860 1260
rect 2920 1180 3060 1260
rect 930 1170 990 1180
rect 1480 1170 1540 1180
rect 2310 1170 2370 1180
rect 2860 1170 2920 1180
rect 3420 1020 3660 1800
rect 580 980 660 990
rect 1120 980 1180 990
rect 1660 980 1720 990
rect 2120 980 2180 990
rect 2680 980 2740 990
rect 560 900 580 980
rect 660 900 1120 980
rect 1180 900 1660 980
rect 1720 900 2120 980
rect 2180 900 2680 980
rect 2740 900 3060 980
rect 3420 950 3940 1020
rect 580 890 660 900
rect 1120 890 1180 900
rect 1660 890 1720 900
rect 2120 890 2180 900
rect 2680 890 2740 900
rect 3420 830 3480 950
rect 3540 830 3810 950
rect 3870 830 3940 950
rect 140 820 220 830
rect 1020 820 1080 830
rect 1570 820 1630 830
rect 2210 820 2270 830
rect 2770 820 2830 830
rect 3420 820 3940 830
rect 80 740 140 820
rect 220 740 1020 820
rect 1080 740 1570 820
rect 1630 740 2210 820
rect 2270 740 2770 820
rect 2830 740 3060 820
rect 140 730 220 740
rect 1020 730 1080 740
rect 1570 730 1630 740
rect 2210 730 2270 740
rect 2770 730 2830 740
rect 3640 650 3700 660
rect 3320 640 3380 650
rect 3110 630 3200 640
rect 280 590 360 600
rect 280 430 290 590
rect 350 430 360 590
rect 3080 550 3110 630
rect 3200 550 3320 630
rect 3380 550 3640 630
rect 3110 540 3200 550
rect 3320 540 3380 550
rect 280 400 360 430
rect 840 440 920 450
rect 280 300 840 400
rect 900 400 920 440
rect 1280 440 1460 450
rect 1280 400 1300 440
rect 900 300 1300 400
rect 900 280 920 300
rect 840 270 920 280
rect 1280 280 1300 300
rect 1440 400 1460 440
rect 1840 440 2020 450
rect 1440 300 1840 400
rect 1440 280 1460 300
rect 1280 270 1460 280
rect 2000 400 2020 440
rect 2400 440 2580 450
rect 2000 300 2400 400
rect 2000 280 2020 300
rect 1840 270 2020 280
rect 2550 400 2580 440
rect 2920 440 3010 450
rect 2920 400 2950 440
rect 2550 300 2950 400
rect 2550 280 2580 300
rect 2400 270 2580 280
rect 2920 280 2950 300
rect 3980 640 4040 650
rect 3700 550 3980 630
rect 4090 640 4150 650
rect 4040 550 4090 630
rect 4150 550 4180 630
rect 3980 540 4040 550
rect 4090 540 4150 550
rect 3640 430 3700 440
rect 2920 270 3010 280
rect -40 180 3960 190
rect -40 120 200 180
rect 270 120 360 180
rect 430 120 3400 180
rect 3470 120 3560 180
rect 3630 120 3720 180
rect 3790 120 3880 180
rect 3950 120 3960 180
rect -40 110 170 120
rect 200 110 270 120
rect 360 110 430 120
rect 3400 110 3470 120
rect 3560 110 3630 120
rect 3720 110 3790 120
rect 3880 110 3950 120
<< via2 >>
rect 2980 2740 3080 2960
rect 1660 1860 1670 1980
rect 1670 1860 1730 1980
rect 1730 1860 1740 1980
rect 4140 1880 4320 2040
rect 940 1520 1060 1620
<< metal3 >>
rect 2970 2960 3090 2965
rect 2970 2740 2980 2960
rect 3080 2740 3220 2960
rect 2970 2735 3090 2740
rect 4130 2040 4330 2045
rect 560 1980 1760 2000
rect 560 1860 1660 1980
rect 1740 1860 1760 1980
rect 4130 1880 4140 2040
rect 4320 1880 4330 2040
rect 4130 1875 4330 1880
rect 560 1840 1760 1860
rect 930 1620 1070 1625
rect 870 1480 880 1620
rect 1120 1480 1130 1620
<< via3 >>
rect 4140 1880 4320 2040
rect 880 1520 940 1620
rect 940 1520 1060 1620
rect 1060 1520 1120 1620
rect 880 1480 1120 1520
<< metal4 >>
rect 4139 2040 4321 2041
rect 160 1600 320 1920
rect 3740 1880 4140 2040
rect 4320 1880 4360 2040
rect 4139 1879 4321 1880
rect 940 1680 1060 1720
rect 840 1621 1120 1680
rect 840 1620 1121 1621
rect 840 1600 880 1620
rect 160 1480 880 1600
rect 1120 1480 1121 1620
rect 160 1479 1121 1480
rect 160 1440 1120 1479
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_0
timestamp 1762739948
transform 1 0 386 0 1 1960
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_K8PL49  sky130_fd_pr__cap_mim_m3_1_K8PL49_0
timestamp 1762739948
transform 0 -1 3500 1 0 2386
box -586 -440 586 440
use sky130_fd_pr__nfet_03v3_nvt_7WRH84  sky130_fd_pr__nfet_03v3_nvt_7WRH84_0
timestamp 1762739948
transform 1 0 1924 0 1 618
box -1244 -658 1244 658
use sky130_fd_pr__nfet_g5v0d10v5_HU3XD6  sky130_fd_pr__nfet_g5v0d10v5_HU3XD6_0
timestamp 1762739948
transform 1 0 317 0 1 418
box -357 -458 357 458
use sky130_fd_pr__nfet_g5v0d10v5_R4FM4P  sky130_fd_pr__nfet_g5v0d10v5_R4FM4P_0
timestamp 1762739948
transform 1 0 3675 0 1 618
box -515 -658 515 658
use sky130_fd_pr__pfet_g5v0d10v5_F6REXY  sky130_fd_pr__pfet_g5v0d10v5_F6REXY_0
timestamp 1762739948
transform 1 0 -713 0 1 1937
box -447 -497 447 497
use sky130_fd_pr__pfet_g5v0d10v5_ZPAR4F  sky130_fd_pr__pfet_g5v0d10v5_ZPAR4F_0
timestamp 1762739948
transform 1 0 2021 0 1 2137
box -861 -697 861 697
<< labels >>
flabel metal2 -40 1180 40 1260 0 FreeSans 960 0 0 0 IN_N
port 0 nsew
flabel metal2 -40 1340 40 1420 0 FreeSans 960 0 0 0 IN_P
port 1 nsew
flabel metal1 140 940 220 1000 0 FreeSans 640 0 0 0 VN
flabel metal2 3420 1420 3660 1690 0 FreeSans 640 0 0 0 VOUT
port 2 nsew
flabel metal1 100 2600 380 2840 0 FreeSans 960 0 0 0 VDD
port 3 nsew
flabel metal1 80 -240 360 0 0 FreeSans 960 0 0 0 VSS
port 4 nsew
flabel metal2 -40 110 40 190 0 FreeSans 960 0 0 0 VBIASN_G5W2L1
port 5 nsew
flabel metal1 860 1600 940 1680 0 FreeSans 640 0 0 0 VOUTSTAGE1
<< end >>
