magic
tech sky130A
magscale 1 2
timestamp 1762739948
<< pwell >>
rect -278 -658 278 658
<< mvnmos >>
rect -50 -400 50 400
<< mvndiff >>
rect -108 388 -50 400
rect -108 -388 -96 388
rect -62 -388 -50 388
rect -108 -400 -50 -388
rect 50 388 108 400
rect 50 -388 62 388
rect 96 -388 108 388
rect 50 -400 108 -388
<< mvndiffc >>
rect -96 -388 -62 388
rect 62 -388 96 388
<< mvpsubdiff >>
rect -242 610 242 622
rect -242 576 -134 610
rect 134 576 242 610
rect -242 564 242 576
rect -242 514 -184 564
rect -242 -514 -230 514
rect -196 -514 -184 514
rect 184 514 242 564
rect -242 -564 -184 -514
rect 184 -514 196 514
rect 230 -514 242 514
rect 184 -564 242 -514
rect -242 -576 242 -564
rect -242 -610 -134 -576
rect 134 -610 242 -576
rect -242 -622 242 -610
<< mvpsubdiffcont >>
rect -134 576 134 610
rect -230 -514 -196 514
rect 196 -514 230 514
rect -134 -610 134 -576
<< poly >>
rect -50 472 50 488
rect -50 438 -34 472
rect 34 438 50 472
rect -50 400 50 438
rect -50 -438 50 -400
rect -50 -472 -34 -438
rect 34 -472 50 -438
rect -50 -488 50 -472
<< polycont >>
rect -34 438 34 472
rect -34 -472 34 -438
<< locali >>
rect -230 576 -134 610
rect 134 576 230 610
rect -230 514 -196 576
rect 196 514 230 576
rect -50 438 -34 472
rect 34 438 50 472
rect -96 388 -62 404
rect -96 -404 -62 -388
rect 62 388 96 404
rect 62 -404 96 -388
rect -50 -472 -34 -438
rect 34 -472 50 -438
rect -230 -576 -196 -514
rect 196 -576 230 -514
rect -230 -610 -134 -576
rect 134 -610 230 -576
<< viali >>
rect -34 438 34 472
rect -230 -230 -196 230
rect -96 -155 -62 155
rect 62 61 96 371
rect 196 -230 230 230
rect -34 -472 34 -438
rect -78 -610 78 -576
<< metal1 >>
rect -46 472 46 478
rect -46 438 -34 472
rect 34 438 46 472
rect -46 432 46 438
rect 56 371 102 383
rect -236 230 -190 242
rect -236 -230 -230 230
rect -196 -230 -190 230
rect -102 155 -56 167
rect -102 -155 -96 155
rect -62 -155 -56 155
rect 56 61 62 371
rect 96 61 102 371
rect 56 49 102 61
rect 190 230 236 242
rect -102 -167 -56 -155
rect -236 -242 -190 -230
rect 190 -230 196 230
rect 230 -230 236 230
rect 190 -242 236 -230
rect -46 -438 46 -432
rect -46 -472 -34 -438
rect 34 -472 46 -438
rect -46 -478 46 -472
rect -90 -576 90 -570
rect -90 -610 -78 -576
rect 78 -610 90 -576
rect -90 -616 90 -610
<< properties >>
string FIXED_BBOX -213 -593 213 593
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -40 viadrn 40 viagate 100 viagb 40 viagr 40 viagl 40 viagt 0
<< end >>
