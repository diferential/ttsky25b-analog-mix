magic
tech sky130A
magscale 1 2
timestamp 1720441783
<< error_p >>
rect -29 132 29 138
rect -29 98 -17 132
rect -29 92 29 98
rect -29 -98 29 -92
rect -29 -132 -17 -98
rect -29 -138 29 -132
<< pwell >>
rect -226 -270 226 270
<< nmos >>
rect -30 -60 30 60
<< ndiff >>
rect -88 48 -30 60
rect -88 -48 -76 48
rect -42 -48 -30 48
rect -88 -60 -30 -48
rect 30 48 88 60
rect 30 -48 42 48
rect 76 -48 88 48
rect 30 -60 88 -48
<< ndiffc >>
rect -76 -48 -42 48
rect 42 -48 76 48
<< psubdiff >>
rect -190 200 190 234
rect -190 -200 -156 200
rect 156 -200 190 200
rect -190 -234 -94 -200
rect 94 -234 190 -200
<< psubdiffcont >>
rect -94 -234 94 -200
<< poly >>
rect -33 132 33 148
rect -33 98 -17 132
rect 17 98 33 132
rect -33 82 33 98
rect -30 60 30 82
rect -30 -82 30 -60
rect -33 -98 33 -82
rect -33 -132 -17 -98
rect 17 -132 33 -98
rect -33 -148 33 -132
<< polycont >>
rect -17 98 17 132
rect -17 -132 17 -98
<< locali >>
rect -33 98 -17 132
rect 17 98 33 132
rect -76 48 -42 64
rect -76 -64 -42 -48
rect 42 48 76 64
rect 42 -64 76 -48
rect -33 -132 -17 -98
rect 17 -132 33 -98
rect -110 -234 -94 -200
rect 94 -234 110 -200
<< viali >>
rect -17 98 17 132
rect -76 -48 -42 48
rect 42 -48 76 48
rect -17 -132 17 -98
<< metal1 >>
rect -29 132 29 138
rect -29 98 -17 132
rect 17 98 29 132
rect -29 92 29 98
rect -82 48 -36 60
rect -82 -48 -76 48
rect -42 -48 -36 48
rect -82 -60 -36 -48
rect 36 48 82 60
rect 36 -48 42 48
rect 76 -48 82 48
rect 36 -60 82 -48
rect -29 -98 29 -92
rect -29 -132 -17 -98
rect 17 -132 29 -98
rect -29 -138 29 -132
<< properties >>
string FIXED_BBOX -173 -217 173 217
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.600 l 0.300 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
