magic
tech sky130A
magscale 1 2
timestamp 1724417029
<< nwell >>
rect -387 -497 387 497
<< mvpmos >>
rect -129 -200 -29 200
rect 29 -200 129 200
<< mvpdiff >>
rect -187 188 -129 200
rect -187 -188 -175 188
rect -141 -188 -129 188
rect -187 -200 -129 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 129 188 187 200
rect 129 -188 141 188
rect 175 -188 187 188
rect 129 -200 187 -188
<< mvpdiffc >>
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
<< mvnsubdiff >>
rect -321 419 321 431
rect -321 385 -213 419
rect 213 385 321 419
rect -321 373 321 385
rect -321 323 -263 373
rect -321 -323 -309 323
rect -275 -323 -263 323
rect 263 323 321 373
rect -321 -373 -263 -323
rect 263 -323 275 323
rect 309 -323 321 323
rect 263 -373 321 -323
rect -321 -385 321 -373
rect -321 -419 -213 -385
rect 213 -419 321 -385
rect -321 -431 321 -419
<< mvnsubdiffcont >>
rect -213 385 213 419
rect -309 -323 -275 323
rect 275 -323 309 323
rect -213 -419 213 -385
<< poly >>
rect -129 281 -29 297
rect -129 247 -113 281
rect -45 247 -29 281
rect -129 200 -29 247
rect 29 281 129 297
rect 29 247 45 281
rect 113 247 129 281
rect 29 200 129 247
rect -129 -247 -29 -200
rect -129 -281 -113 -247
rect -45 -281 -29 -247
rect -129 -297 -29 -281
rect 29 -247 129 -200
rect 29 -281 45 -247
rect 113 -281 129 -247
rect 29 -297 129 -281
<< polycont >>
rect -113 247 -45 281
rect 45 247 113 281
rect -113 -281 -45 -247
rect 45 -281 113 -247
<< locali >>
rect -309 385 -213 419
rect 213 385 309 419
rect -309 323 -275 385
rect 275 323 309 385
rect -129 247 -113 281
rect -45 247 -29 281
rect 29 247 45 281
rect 113 247 129 281
rect -175 188 -141 204
rect -175 -204 -141 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 141 188 175 204
rect 141 -204 175 -188
rect -129 -281 -113 -247
rect -45 -281 -29 -247
rect 29 -281 45 -247
rect 113 -281 129 -247
rect -309 -385 -275 -323
rect 275 -385 309 -323
rect -309 -419 -213 -385
rect 213 -419 309 -385
<< viali >>
rect -113 247 -45 281
rect 45 247 113 281
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect -113 -281 -45 -247
rect 45 -281 113 -247
rect -138 -419 138 -385
<< metal1 >>
rect -125 281 -33 287
rect -125 247 -113 281
rect -45 247 -33 281
rect -125 241 -33 247
rect 33 281 125 287
rect 33 247 45 281
rect 113 247 125 281
rect 33 241 125 247
rect -181 188 -135 200
rect -181 -188 -175 188
rect -141 -188 -135 188
rect -181 -200 -135 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 135 188 181 200
rect 135 -188 141 188
rect 175 -188 181 188
rect 135 -200 181 -188
rect -125 -247 -33 -241
rect -125 -281 -113 -247
rect -45 -281 -33 -247
rect -125 -287 -33 -281
rect 33 -247 125 -241
rect 33 -281 45 -247
rect 113 -281 125 -247
rect 33 -287 125 -281
rect -150 -385 150 -379
rect -150 -419 -138 -385
rect 138 -419 150 -385
rect -150 -425 150 -419
<< properties >>
string FIXED_BBOX -292 -402 292 402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 50 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__pfet_g5v0d10v5_3827BU gencell
<< end >>
