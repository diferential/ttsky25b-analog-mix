magic
tech sky130A
magscale 1 2
timestamp 1725637093
<< error_p >>
rect -31 -111 31 -105
rect -31 -145 -19 -111
rect -31 -151 31 -145
<< nwell >>
rect -231 -284 231 284
<< pmoslvt >>
rect -35 -64 35 136
<< pdiff >>
rect -93 124 -35 136
rect -93 -52 -81 124
rect -47 -52 -35 124
rect -93 -64 -35 -52
rect 35 124 93 136
rect 35 -52 47 124
rect 81 -52 93 124
rect 35 -64 93 -52
<< pdiffc >>
rect -81 -52 -47 124
rect 47 -52 81 124
<< nsubdiff >>
rect -195 214 195 248
rect -195 151 -161 214
rect 161 151 195 214
rect -195 -214 -161 -151
rect 161 -214 195 -151
rect -195 -248 -99 -214
rect 99 -248 195 -214
<< nsubdiffcont >>
rect -195 -151 -161 151
rect 161 -151 195 151
rect -99 -248 99 -214
<< poly >>
rect -35 136 35 162
rect -35 -111 35 -64
rect -35 -145 -19 -111
rect 19 -145 35 -111
rect -35 -161 35 -145
<< polycont >>
rect -19 -145 19 -111
<< locali >>
rect -195 151 -161 248
rect 161 151 195 248
rect -81 124 -47 140
rect -81 -68 -47 -52
rect 47 124 81 140
rect 47 -68 81 -52
rect -35 -145 -19 -111
rect 19 -145 35 -111
rect -195 -214 -161 -151
rect 161 -214 195 -151
rect -195 -248 -99 -214
rect 99 -248 195 -214
<< viali >>
rect -161 214 161 248
rect -81 -52 -47 124
rect 47 -52 81 124
rect -19 -145 19 -111
<< metal1 >>
rect -173 248 173 254
rect -173 214 -161 248
rect 161 214 173 248
rect -173 208 173 214
rect -87 124 -41 136
rect -87 -52 -81 124
rect -47 -52 -41 124
rect -87 -64 -41 -52
rect 41 124 87 136
rect 41 -52 47 124
rect 81 -52 87 124
rect 41 -64 87 -52
rect -31 -111 31 -105
rect -31 -145 -19 -111
rect 19 -145 31 -111
rect -31 -151 31 -145
<< properties >>
string FIXED_BBOX -178 -231 178 231
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 100
<< end >>
