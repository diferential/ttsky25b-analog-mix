magic
tech sky130A
magscale 1 2
timestamp 1725323004
<< pwell >>
rect -278 -4221 278 4221
<< nnmos >>
rect -50 3163 50 3963
rect -50 2145 50 2945
rect -50 1127 50 1927
rect -50 109 50 909
rect -50 -909 50 -109
rect -50 -1927 50 -1127
rect -50 -2945 50 -2145
rect -50 -3963 50 -3163
<< mvndiff >>
rect -108 3951 -50 3963
rect -108 3175 -96 3951
rect -62 3175 -50 3951
rect -108 3163 -50 3175
rect 50 3951 108 3963
rect 50 3175 62 3951
rect 96 3175 108 3951
rect 50 3163 108 3175
rect -108 2933 -50 2945
rect -108 2157 -96 2933
rect -62 2157 -50 2933
rect -108 2145 -50 2157
rect 50 2933 108 2945
rect 50 2157 62 2933
rect 96 2157 108 2933
rect 50 2145 108 2157
rect -108 1915 -50 1927
rect -108 1139 -96 1915
rect -62 1139 -50 1915
rect -108 1127 -50 1139
rect 50 1915 108 1927
rect 50 1139 62 1915
rect 96 1139 108 1915
rect 50 1127 108 1139
rect -108 897 -50 909
rect -108 121 -96 897
rect -62 121 -50 897
rect -108 109 -50 121
rect 50 897 108 909
rect 50 121 62 897
rect 96 121 108 897
rect 50 109 108 121
rect -108 -121 -50 -109
rect -108 -897 -96 -121
rect -62 -897 -50 -121
rect -108 -909 -50 -897
rect 50 -121 108 -109
rect 50 -897 62 -121
rect 96 -897 108 -121
rect 50 -909 108 -897
rect -108 -1139 -50 -1127
rect -108 -1915 -96 -1139
rect -62 -1915 -50 -1139
rect -108 -1927 -50 -1915
rect 50 -1139 108 -1127
rect 50 -1915 62 -1139
rect 96 -1915 108 -1139
rect 50 -1927 108 -1915
rect -108 -2157 -50 -2145
rect -108 -2933 -96 -2157
rect -62 -2933 -50 -2157
rect -108 -2945 -50 -2933
rect 50 -2157 108 -2145
rect 50 -2933 62 -2157
rect 96 -2933 108 -2157
rect 50 -2945 108 -2933
rect -108 -3175 -50 -3163
rect -108 -3951 -96 -3175
rect -62 -3951 -50 -3175
rect -108 -3963 -50 -3951
rect 50 -3175 108 -3163
rect 50 -3951 62 -3175
rect 96 -3951 108 -3175
rect 50 -3963 108 -3951
<< mvndiffc >>
rect -96 3175 -62 3951
rect 62 3175 96 3951
rect -96 2157 -62 2933
rect 62 2157 96 2933
rect -96 1139 -62 1915
rect 62 1139 96 1915
rect -96 121 -62 897
rect 62 121 96 897
rect -96 -897 -62 -121
rect 62 -897 96 -121
rect -96 -1915 -62 -1139
rect 62 -1915 96 -1139
rect -96 -2933 -62 -2157
rect 62 -2933 96 -2157
rect -96 -3951 -62 -3175
rect 62 -3951 96 -3175
<< mvpsubdiff >>
rect -242 4173 242 4185
rect -242 4139 -134 4173
rect 134 4139 242 4173
rect -242 4127 242 4139
rect -242 4077 -184 4127
rect -242 -4077 -230 4077
rect -196 -4077 -184 4077
rect 184 4077 242 4127
rect -242 -4127 -184 -4077
rect 184 -4077 196 4077
rect 230 -4077 242 4077
rect 184 -4127 242 -4077
rect -242 -4139 242 -4127
rect -242 -4173 -134 -4139
rect 134 -4173 242 -4139
rect -242 -4185 242 -4173
<< mvpsubdiffcont >>
rect -134 4139 134 4173
rect -230 -4077 -196 4077
rect 196 -4077 230 4077
rect -134 -4173 134 -4139
<< poly >>
rect -50 4035 50 4051
rect -50 4001 -34 4035
rect 34 4001 50 4035
rect -50 3963 50 4001
rect -50 3125 50 3163
rect -50 3091 -34 3125
rect 34 3091 50 3125
rect -50 3075 50 3091
rect -50 3017 50 3033
rect -50 2983 -34 3017
rect 34 2983 50 3017
rect -50 2945 50 2983
rect -50 2107 50 2145
rect -50 2073 -34 2107
rect 34 2073 50 2107
rect -50 2057 50 2073
rect -50 1999 50 2015
rect -50 1965 -34 1999
rect 34 1965 50 1999
rect -50 1927 50 1965
rect -50 1089 50 1127
rect -50 1055 -34 1089
rect 34 1055 50 1089
rect -50 1039 50 1055
rect -50 981 50 997
rect -50 947 -34 981
rect 34 947 50 981
rect -50 909 50 947
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -947 50 -909
rect -50 -981 -34 -947
rect 34 -981 50 -947
rect -50 -997 50 -981
rect -50 -1055 50 -1039
rect -50 -1089 -34 -1055
rect 34 -1089 50 -1055
rect -50 -1127 50 -1089
rect -50 -1965 50 -1927
rect -50 -1999 -34 -1965
rect 34 -1999 50 -1965
rect -50 -2015 50 -1999
rect -50 -2073 50 -2057
rect -50 -2107 -34 -2073
rect 34 -2107 50 -2073
rect -50 -2145 50 -2107
rect -50 -2983 50 -2945
rect -50 -3017 -34 -2983
rect 34 -3017 50 -2983
rect -50 -3033 50 -3017
rect -50 -3091 50 -3075
rect -50 -3125 -34 -3091
rect 34 -3125 50 -3091
rect -50 -3163 50 -3125
rect -50 -4001 50 -3963
rect -50 -4035 -34 -4001
rect 34 -4035 50 -4001
rect -50 -4051 50 -4035
<< polycont >>
rect -34 4001 34 4035
rect -34 3091 34 3125
rect -34 2983 34 3017
rect -34 2073 34 2107
rect -34 1965 34 1999
rect -34 1055 34 1089
rect -34 947 34 981
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -981 34 -947
rect -34 -1089 34 -1055
rect -34 -1999 34 -1965
rect -34 -2107 34 -2073
rect -34 -3017 34 -2983
rect -34 -3125 34 -3091
rect -34 -4035 34 -4001
<< locali >>
rect -230 4139 -134 4173
rect 134 4139 230 4173
rect -230 4077 -196 4139
rect 196 4077 230 4139
rect -50 4001 -34 4035
rect 34 4001 50 4035
rect -96 3951 -62 3967
rect -96 3159 -62 3175
rect 62 3951 96 3967
rect 62 3159 96 3175
rect -50 3091 -34 3125
rect 34 3091 50 3125
rect -50 2983 -34 3017
rect 34 2983 50 3017
rect -96 2933 -62 2949
rect -96 2141 -62 2157
rect 62 2933 96 2949
rect 62 2141 96 2157
rect -50 2073 -34 2107
rect 34 2073 50 2107
rect -50 1965 -34 1999
rect 34 1965 50 1999
rect -96 1915 -62 1931
rect -96 1123 -62 1139
rect 62 1915 96 1931
rect 62 1123 96 1139
rect -50 1055 -34 1089
rect 34 1055 50 1089
rect -50 947 -34 981
rect 34 947 50 981
rect -96 897 -62 913
rect -96 105 -62 121
rect 62 897 96 913
rect 62 105 96 121
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -913 -62 -897
rect 62 -121 96 -105
rect 62 -913 96 -897
rect -50 -981 -34 -947
rect 34 -981 50 -947
rect -50 -1089 -34 -1055
rect 34 -1089 50 -1055
rect -96 -1139 -62 -1123
rect -96 -1931 -62 -1915
rect 62 -1139 96 -1123
rect 62 -1931 96 -1915
rect -50 -1999 -34 -1965
rect 34 -1999 50 -1965
rect -50 -2107 -34 -2073
rect 34 -2107 50 -2073
rect -96 -2157 -62 -2141
rect -96 -2949 -62 -2933
rect 62 -2157 96 -2141
rect 62 -2949 96 -2933
rect -50 -3017 -34 -2983
rect 34 -3017 50 -2983
rect -50 -3125 -34 -3091
rect 34 -3125 50 -3091
rect -96 -3175 -62 -3159
rect -96 -3967 -62 -3951
rect 62 -3175 96 -3159
rect 62 -3967 96 -3951
rect -50 -4035 -34 -4001
rect 34 -4035 50 -4001
rect -230 -4139 -196 -4077
rect 196 -4139 230 -4077
rect -230 -4173 -134 -4139
rect 134 -4173 230 -4139
<< viali >>
rect -34 4001 34 4035
rect -96 3192 -62 3502
rect 62 3624 96 3934
rect -34 3091 34 3125
rect -34 2983 34 3017
rect -96 2174 -62 2484
rect 62 2606 96 2916
rect -34 2073 34 2107
rect -34 1965 34 1999
rect -96 1156 -62 1466
rect 62 1588 96 1898
rect -34 1055 34 1089
rect -34 947 34 981
rect -96 138 -62 448
rect 62 570 96 880
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -880 -62 -570
rect 62 -448 96 -138
rect -34 -981 34 -947
rect -34 -1089 34 -1055
rect -96 -1898 -62 -1588
rect 62 -1466 96 -1156
rect -34 -1999 34 -1965
rect -34 -2107 34 -2073
rect -96 -2916 -62 -2606
rect 62 -2484 96 -2174
rect -34 -3017 34 -2983
rect -34 -3125 34 -3091
rect -96 -3934 -62 -3624
rect 62 -3502 96 -3192
rect -34 -4035 34 -4001
rect -118 -4173 118 -4139
<< metal1 >>
rect -46 4035 46 4041
rect -46 4001 -34 4035
rect 34 4001 46 4035
rect -46 3995 46 4001
rect 56 3934 102 3946
rect 56 3624 62 3934
rect 96 3624 102 3934
rect 56 3612 102 3624
rect -102 3502 -56 3514
rect -102 3192 -96 3502
rect -62 3192 -56 3502
rect -102 3180 -56 3192
rect -46 3125 46 3131
rect -46 3091 -34 3125
rect 34 3091 46 3125
rect -46 3085 46 3091
rect -46 3017 46 3023
rect -46 2983 -34 3017
rect 34 2983 46 3017
rect -46 2977 46 2983
rect 56 2916 102 2928
rect 56 2606 62 2916
rect 96 2606 102 2916
rect 56 2594 102 2606
rect -102 2484 -56 2496
rect -102 2174 -96 2484
rect -62 2174 -56 2484
rect -102 2162 -56 2174
rect -46 2107 46 2113
rect -46 2073 -34 2107
rect 34 2073 46 2107
rect -46 2067 46 2073
rect -46 1999 46 2005
rect -46 1965 -34 1999
rect 34 1965 46 1999
rect -46 1959 46 1965
rect 56 1898 102 1910
rect 56 1588 62 1898
rect 96 1588 102 1898
rect 56 1576 102 1588
rect -102 1466 -56 1478
rect -102 1156 -96 1466
rect -62 1156 -56 1466
rect -102 1144 -56 1156
rect -46 1089 46 1095
rect -46 1055 -34 1089
rect 34 1055 46 1089
rect -46 1049 46 1055
rect -46 981 46 987
rect -46 947 -34 981
rect 34 947 46 981
rect -46 941 46 947
rect 56 880 102 892
rect 56 570 62 880
rect 96 570 102 880
rect 56 558 102 570
rect -102 448 -56 460
rect -102 138 -96 448
rect -62 138 -56 448
rect -102 126 -56 138
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect 56 -138 102 -126
rect 56 -448 62 -138
rect 96 -448 102 -138
rect 56 -460 102 -448
rect -102 -570 -56 -558
rect -102 -880 -96 -570
rect -62 -880 -56 -570
rect -102 -892 -56 -880
rect -46 -947 46 -941
rect -46 -981 -34 -947
rect 34 -981 46 -947
rect -46 -987 46 -981
rect -46 -1055 46 -1049
rect -46 -1089 -34 -1055
rect 34 -1089 46 -1055
rect -46 -1095 46 -1089
rect 56 -1156 102 -1144
rect 56 -1466 62 -1156
rect 96 -1466 102 -1156
rect 56 -1478 102 -1466
rect -102 -1588 -56 -1576
rect -102 -1898 -96 -1588
rect -62 -1898 -56 -1588
rect -102 -1910 -56 -1898
rect -46 -1965 46 -1959
rect -46 -1999 -34 -1965
rect 34 -1999 46 -1965
rect -46 -2005 46 -1999
rect -46 -2073 46 -2067
rect -46 -2107 -34 -2073
rect 34 -2107 46 -2073
rect -46 -2113 46 -2107
rect 56 -2174 102 -2162
rect 56 -2484 62 -2174
rect 96 -2484 102 -2174
rect 56 -2496 102 -2484
rect -102 -2606 -56 -2594
rect -102 -2916 -96 -2606
rect -62 -2916 -56 -2606
rect -102 -2928 -56 -2916
rect -46 -2983 46 -2977
rect -46 -3017 -34 -2983
rect 34 -3017 46 -2983
rect -46 -3023 46 -3017
rect -46 -3091 46 -3085
rect -46 -3125 -34 -3091
rect 34 -3125 46 -3091
rect -46 -3131 46 -3125
rect 56 -3192 102 -3180
rect 56 -3502 62 -3192
rect 96 -3502 102 -3192
rect 56 -3514 102 -3502
rect -102 -3624 -56 -3612
rect -102 -3934 -96 -3624
rect -62 -3934 -56 -3624
rect -102 -3946 -56 -3934
rect -46 -4001 46 -3995
rect -46 -4035 -34 -4001
rect 34 -4035 46 -4001
rect -46 -4041 46 -4035
rect -130 -4139 130 -4133
rect -130 -4173 -118 -4139
rect 118 -4173 130 -4139
rect -130 -4179 130 -4173
<< properties >>
string FIXED_BBOX -213 -4156 213 4156
string gencell sky130_fd_pr__nfet_03v3_nvt
string library sky130
string parameters w 4 l 0.5 m 8 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -40 viadrn +40 viagate 100 viagb 60 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__nfet_03v3_nvt_7FJT7R gencell
<< end >>
