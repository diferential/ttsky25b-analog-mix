magic
tech sky130A
magscale 1 2
timestamp 1720441783
<< error_p >>
rect -88 -101 -30 -95
rect 30 -101 88 -95
rect -88 -135 -76 -101
rect 30 -135 42 -101
rect -88 -141 -30 -135
rect 30 -141 88 -135
<< nwell >>
rect -285 -274 285 274
<< pmos >>
rect -89 -54 -29 126
rect 29 -54 89 126
<< pdiff >>
rect -147 114 -89 126
rect -147 -42 -135 114
rect -101 -42 -89 114
rect -147 -54 -89 -42
rect -29 114 29 126
rect -29 -42 -17 114
rect 17 -42 29 114
rect -29 -54 29 -42
rect 89 114 147 126
rect 89 -42 101 114
rect 135 -42 147 114
rect 89 -54 147 -42
<< pdiffc >>
rect -135 -42 -101 114
rect -17 -42 17 114
rect 101 -42 135 114
<< nsubdiff >>
rect -249 204 -153 238
rect 153 204 249 238
rect -249 -204 -215 204
rect 215 -204 249 204
rect -249 -238 249 -204
<< nsubdiffcont >>
rect -153 204 153 238
<< poly >>
rect -89 126 -29 152
rect 29 126 89 152
rect -89 -85 -29 -54
rect 29 -85 89 -54
rect -92 -101 -26 -85
rect -92 -135 -76 -101
rect -42 -135 -26 -101
rect -92 -151 -26 -135
rect 26 -101 92 -85
rect 26 -135 42 -101
rect 76 -135 92 -101
rect 26 -151 92 -135
<< polycont >>
rect -76 -135 -42 -101
rect 42 -135 76 -101
<< locali >>
rect -169 204 -153 238
rect 153 204 169 238
rect -135 114 -101 130
rect -135 -58 -101 -42
rect -17 114 17 130
rect -17 -58 17 -42
rect 101 114 135 130
rect 101 -58 135 -42
rect -92 -135 -76 -101
rect -42 -135 -26 -101
rect 26 -135 42 -101
rect 76 -135 92 -101
<< viali >>
rect -135 -42 -101 114
rect -17 -42 17 114
rect 101 -42 135 114
rect -76 -135 -42 -101
rect 42 -135 76 -101
<< metal1 >>
rect -141 114 -95 126
rect -141 -42 -135 114
rect -101 -42 -95 114
rect -141 -54 -95 -42
rect -23 114 23 126
rect -23 -42 -17 114
rect 17 -42 23 114
rect -23 -54 23 -42
rect 95 114 141 126
rect 95 -42 101 114
rect 135 -42 141 114
rect 95 -54 141 -42
rect -88 -101 -30 -95
rect -88 -135 -76 -101
rect -42 -135 -30 -101
rect -88 -141 -30 -135
rect 30 -101 88 -95
rect 30 -135 42 -101
rect 76 -135 88 -101
rect 30 -141 88 -135
<< properties >>
string FIXED_BBOX -232 -221 232 221
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.90 l 0.30 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
