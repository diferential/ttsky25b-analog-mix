magic
tech sky130A
magscale 1 2
timestamp 1720618976
<< nmoslvt >>
rect -25 -50 25 50
<< ndiff >>
rect -83 38 -25 50
rect -83 -38 -71 38
rect -37 -38 -25 38
rect -83 -50 -25 -38
rect 25 38 83 50
rect 25 -38 37 38
rect 71 -38 83 38
rect 25 -50 83 -38
<< ndiffc >>
rect -71 -38 -37 38
rect 37 -38 71 38
<< poly >>
rect -25 50 25 76
rect -25 -76 25 -50
<< locali >>
rect -71 38 -37 54
rect -71 -54 -37 -38
rect 37 38 71 54
rect 37 -54 71 -38
<< viali >>
rect -71 -38 -37 38
rect 37 -38 71 38
<< metal1 >>
rect -77 38 -31 50
rect -77 -38 -71 38
rect -37 -38 -31 38
rect -77 -50 -31 -38
rect 31 38 77 50
rect 31 -38 37 38
rect 71 -38 77 38
rect 31 -50 77 -38
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 0.5 l 0.25 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
